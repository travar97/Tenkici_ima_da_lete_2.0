
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);
	
	port
	(
		clk_i    : in  std_logic;
		addr_i	: in  unsigned( ADDR_WIDTH-1 downto 0 );
		data_o	: out	std_logic_vector( DATA_WIDTH-1 downto 0 )
	);
end entity ram;

architecture arch of ram is

	type	ram_t is array ( 0 to 2**ADDR_WIDTH-1 ) of std_logic_vector( DATA_WIDTH-1 downto 0 );
	
-- GENERATED BY BC_MEM_PACKER
-- DATE: Tue Jun 09 11:28:59 2015

	signal mem : ram_t := (


--			***** COLOR PALLETE *****


		0 =>	x"00000080", -- R: 128 G: 0 B: 0
		1 =>	x"00806060", -- R: 96 G: 96 B: 128
		2 =>	x"000040A0", -- R: 160 G: 64 B: 0
		3 =>	x"00000000", -- R: 0 G: 0 B: 0
		4 =>	x"00A4A0A0", -- R: 160 G: 160 B: 164
		5 =>	x"00006000", -- R: 0 G: 96 B: 0
		6 =>	x"00004000", -- R: 0 G: 64 B: 0
		7 =>	x"0000E080", -- R: 128 G: 224 B: 0
		8 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		9 =>	x"00C3C3C3", -- R: 195 G: 195 B: 195
		10 =>	x"00C04040", -- R: 64 G: 64 B: 192
		11 =>	x"00F0CAA6", -- R: 166 G: 202 B: 240
		12 =>	x"00404000", -- R: 0 G: 64 B: 64
		13 =>	x"00800060", -- R: 96 G: 0 B: 128
		14 =>	x"004040C0", -- R: 192 G: 64 B: 64
		15 =>	x"0080E0E0", -- R: 224 G: 224 B: 128
		16 =>	x"0040A0E0", -- R: 224 G: 160 B: 64
		17 =>	x"00006060", -- R: 96 G: 96 B: 0
		18 =>	x"00000000", -- Unused
		19 =>	x"00000000", -- Unused
		20 =>	x"00000000", -- Unused
		21 =>	x"00000000", -- Unused
		22 =>	x"00000000", -- Unused
		23 =>	x"00000000", -- Unused
		24 =>	x"00000000", -- Unused
		25 =>	x"00000000", -- Unused
		26 =>	x"00000000", -- Unused
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused


--			***** 8x8 IMAGES *****


		256 =>	x"00000000", -- IMG_8x8_BRICK
		257 =>	x"01000000",
		258 =>	x"02020202",
		259 =>	x"01000202",
		260 =>	x"02020202",
		261 =>	x"01000202",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01000000",
		265 =>	x"00000000",
		266 =>	x"01000202",
		267 =>	x"02020202",
		268 =>	x"01000202",
		269 =>	x"02020202",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"03030303", -- IMG_8x8_BULLET
		273 =>	x"03030303",
		274 =>	x"03030303",
		275 =>	x"03030303",
		276 =>	x"03030304",
		277 =>	x"03030303",
		278 =>	x"03030404",
		279 =>	x"04030303",
		280 =>	x"03030404",
		281 =>	x"04030303",
		282 =>	x"03030404",
		283 =>	x"04030303",
		284 =>	x"03030303",
		285 =>	x"03030303",
		286 =>	x"03030303",
		287 =>	x"03030303",
		288 =>	x"03050505", -- IMG_8x8_GRASS
		289 =>	x"06050703",
		290 =>	x"05050607",
		291 =>	x"05070507",
		292 =>	x"05050505",
		293 =>	x"05070707",
		294 =>	x"06050507",
		295 =>	x"07060507",
		296 =>	x"05050706",
		297 =>	x"07070706",
		298 =>	x"05060507",
		299 =>	x"07070707",
		300 =>	x"07070707",
		301 =>	x"07060707",
		302 =>	x"03070706",
		303 =>	x"07070703",
		304 =>	x"01040408", -- IMG_8x8_ICE
		305 =>	x"01040408",
		306 =>	x"04040404",
		307 =>	x"04040801",
		308 =>	x"04040404",
		309 =>	x"04080104",
		310 =>	x"08040404",
		311 =>	x"08010404",
		312 =>	x"01040408",
		313 =>	x"01040408",
		314 =>	x"04040801",
		315 =>	x"04040801",
		316 =>	x"04080104",
		317 =>	x"04080104",
		318 =>	x"08010404",
		319 =>	x"08010404",
		320 =>	x"04040404", -- IMG_8x8_IRON
		321 =>	x"04040404",
		322 =>	x"04040404",
		323 =>	x"04040401",
		324 =>	x"04040808",
		325 =>	x"08080101",
		326 =>	x"04040808",
		327 =>	x"08080101",
		328 =>	x"04040808",
		329 =>	x"08080101",
		330 =>	x"04040808",
		331 =>	x"08080101",
		332 =>	x"04040101",
		333 =>	x"01010101",
		334 =>	x"04010101",
		335 =>	x"01010101",
		336 =>	x"01010102", -- IMG_8x8_LIVES_REMAINING_ICON
		337 =>	x"02020101",
		338 =>	x"01020101",
		339 =>	x"02010102",
		340 =>	x"01020102",
		341 =>	x"02020102",
		342 =>	x"01020202",
		343 =>	x"01020202",
		344 =>	x"01020201",
		345 =>	x"01010202",
		346 =>	x"01020202",
		347 =>	x"01020202",
		348 =>	x"01020102",
		349 =>	x"02020102",
		350 =>	x"01020101",
		351 =>	x"02010102",
		352 =>	x"09090909", -- IMG_8x8_NULL
		353 =>	x"09090909",
		354 =>	x"09090909",
		355 =>	x"09090909",
		356 =>	x"09090909",
		357 =>	x"09090909",
		358 =>	x"09090909",
		359 =>	x"09090909",
		360 =>	x"09090909",
		361 =>	x"09090909",
		362 =>	x"09090909",
		363 =>	x"09090909",
		364 =>	x"09090909",
		365 =>	x"09090909",
		366 =>	x"09090909",
		367 =>	x"09090909",
		368 =>	x"01010101", -- IMG_8x8_TANKS_REMAINING_ICON
		369 =>	x"01010101",
		370 =>	x"01030101",
		371 =>	x"03010103",
		372 =>	x"01030103",
		373 =>	x"03030103",
		374 =>	x"01030303",
		375 =>	x"00030303",
		376 =>	x"01030303",
		377 =>	x"00030303",
		378 =>	x"01030103",
		379 =>	x"03030103",
		380 =>	x"01030101",
		381 =>	x"03010103",
		382 =>	x"01010103",
		383 =>	x"03030101",
		384 =>	x"0A0A0A0A", -- IMG_8x8_WATER
		385 =>	x"0A0A0A0B",
		386 =>	x"0A0B0A0A",
		387 =>	x"0A0A0A0A",
		388 =>	x"0A0A0B0A",
		389 =>	x"0A0A0A0A",
		390 =>	x"0A0A0A0B",
		391 =>	x"0A0A0B0A",
		392 =>	x"0A0A0A0A",
		393 =>	x"0A0A0A0B",
		394 =>	x"0A0A0A0B",
		395 =>	x"0A0A0A0A",
		396 =>	x"0A0A0B0A",
		397 =>	x"0B0A0A0A",
		398 =>	x"0B0A0A0A",
		399 =>	x"0A0A0A0A",


--			***** 16x16 IMAGES *****


		400 =>	x"03030303", -- IMG_16x16_BASE_ALIVE
		401 =>	x"03030303",
		402 =>	x"03030303",
		403 =>	x"03030303",
		404 =>	x"01010303",
		405 =>	x"03030303",
		406 =>	x"03030303",
		407 =>	x"03030101",
		408 =>	x"03010103",
		409 =>	x"03030101",
		410 =>	x"01030303",
		411 =>	x"03010103",
		412 =>	x"01010101",
		413 =>	x"03030301",
		414 =>	x"00010303",
		415 =>	x"01010101",
		416 =>	x"03010101",
		417 =>	x"03030301",
		418 =>	x"01030303",
		419 =>	x"01010103",
		420 =>	x"01010101",
		421 =>	x"01010301",
		422 =>	x"01030101",
		423 =>	x"01010101",
		424 =>	x"03030100",
		425 =>	x"01010101",
		426 =>	x"01010101",
		427 =>	x"00010303",
		428 =>	x"03010101",
		429 =>	x"00010101",
		430 =>	x"01010100",
		431 =>	x"01010103",
		432 =>	x"03030101",
		433 =>	x"01010001",
		434 =>	x"01000101",
		435 =>	x"01010303",
		436 =>	x"03030101",
		437 =>	x"01010101",
		438 =>	x"01010101",
		439 =>	x"01010303",
		440 =>	x"03030301",
		441 =>	x"01010301",
		442 =>	x"01030101",
		443 =>	x"01030303",
		444 =>	x"03030303",
		445 =>	x"03030301",
		446 =>	x"01030303",
		447 =>	x"03030303",
		448 =>	x"03030303",
		449 =>	x"03030101",
		450 =>	x"01010303",
		451 =>	x"03030303",
		452 =>	x"03030303",
		453 =>	x"01010101",
		454 =>	x"01010101",
		455 =>	x"03030303",
		456 =>	x"03030303",
		457 =>	x"01010301",
		458 =>	x"01030101",
		459 =>	x"03030303",
		460 =>	x"03030303",
		461 =>	x"03030303",
		462 =>	x"03030303",
		463 =>	x"03030303",
		464 =>	x"03030303", -- IMG_16x16_BASE_DEAD
		465 =>	x"03030303",
		466 =>	x"03030303",
		467 =>	x"03030303",
		468 =>	x"03030303",
		469 =>	x"03020303",
		470 =>	x"03030303",
		471 =>	x"03030303",
		472 =>	x"03030303",
		473 =>	x"02020301",
		474 =>	x"03030303",
		475 =>	x"03030303",
		476 =>	x"03030303",
		477 =>	x"02030101",
		478 =>	x"01030303",
		479 =>	x"03030303",
		480 =>	x"03030302",
		481 =>	x"03010101",
		482 =>	x"01010303",
		483 =>	x"03030303",
		484 =>	x"03030202",
		485 =>	x"03010101",
		486 =>	x"01010101",
		487 =>	x"01030303",
		488 =>	x"03030203",
		489 =>	x"01010101",
		490 =>	x"01010101",
		491 =>	x"01010303",
		492 =>	x"03020203",
		493 =>	x"01010101",
		494 =>	x"01010101",
		495 =>	x"01010303",
		496 =>	x"03020303",
		497 =>	x"01010101",
		498 =>	x"01010101",
		499 =>	x"03010103",
		500 =>	x"03020301",
		501 =>	x"01010101",
		502 =>	x"01030301",
		503 =>	x"03010103",
		504 =>	x"03020303",
		505 =>	x"03010101",
		506 =>	x"03030303",
		507 =>	x"03010303",
		508 =>	x"03020303",
		509 =>	x"03030301",
		510 =>	x"03030303",
		511 =>	x"03010303",
		512 =>	x"03020303",
		513 =>	x"03030303",
		514 =>	x"03030303",
		515 =>	x"03030303",
		516 =>	x"03020303",
		517 =>	x"03030303",
		518 =>	x"03030303",
		519 =>	x"03030303",
		520 =>	x"03020303",
		521 =>	x"03030303",
		522 =>	x"03030303",
		523 =>	x"03030303",
		524 =>	x"03030303",
		525 =>	x"03030303",
		526 =>	x"03030303",
		527 =>	x"03030303",
		528 =>	x"03030303", -- IMG_16x16_BONUS_BOMB
		529 =>	x"03030303",
		530 =>	x"03030303",
		531 =>	x"03030303",
		532 =>	x"03080808",
		533 =>	x"08080808",
		534 =>	x"08080808",
		535 =>	x"08080403",
		536 =>	x"08030303",
		537 =>	x"03030303",
		538 =>	x"03030303",
		539 =>	x"0303080C",
		540 =>	x"08030C0C",
		541 =>	x"0C080808",
		542 =>	x"0404030C",
		543 =>	x"0C0C080C",
		544 =>	x"08030C0C",
		545 =>	x"0C08040C",
		546 =>	x"03030403",
		547 =>	x"0C0C080C",
		548 =>	x"08030C0C",
		549 =>	x"08040404",
		550 =>	x"0C030304",
		551 =>	x"030C080C",
		552 =>	x"08030C08",
		553 =>	x"040C0804",
		554 =>	x"0C040304",
		555 =>	x"030C080C",
		556 =>	x"08030C04",
		557 =>	x"03040303",
		558 =>	x"04030304",
		559 =>	x"030C080C",
		560 =>	x"08030C08",
		561 =>	x"040C0804",
		562 =>	x"0C040304",
		563 =>	x"030C080C",
		564 =>	x"08030C04",
		565 =>	x"03040303",
		566 =>	x"04030304",
		567 =>	x"030C080C",
		568 =>	x"08030C08",
		569 =>	x"040C0804",
		570 =>	x"0C040303",
		571 =>	x"0C0C080C",
		572 =>	x"08030C0C",
		573 =>	x"040C0303",
		574 =>	x"04030C0C",
		575 =>	x"0C0C080C",
		576 =>	x"08030C0C",
		577 =>	x"0C080404",
		578 =>	x"030C0C0C",
		579 =>	x"0C0C080C",
		580 =>	x"08030C0C",
		581 =>	x"0C030303",
		582 =>	x"0C0C0C0C",
		583 =>	x"0C0C080C",
		584 =>	x"04080808",
		585 =>	x"08080808",
		586 =>	x"08080808",
		587 =>	x"0808040C",
		588 =>	x"030C0C0C",
		589 =>	x"0C0C0C0C",
		590 =>	x"0C0C0C0C",
		591 =>	x"0C0C0C03",
		592 =>	x"03030303", -- IMG_16x16_BONUS_GUN
		593 =>	x"03030303",
		594 =>	x"03030303",
		595 =>	x"03030303",
		596 =>	x"03080808",
		597 =>	x"08080808",
		598 =>	x"08080808",
		599 =>	x"08080403",
		600 =>	x"08030303",
		601 =>	x"03030303",
		602 =>	x"03030303",
		603 =>	x"0303080C",
		604 =>	x"08030C0C",
		605 =>	x"0C0C0C0C",
		606 =>	x"0C0C0C0C",
		607 =>	x"0C0C080C",
		608 =>	x"08030C08",
		609 =>	x"0C0C0C0C",
		610 =>	x"0C0C0C0C",
		611 =>	x"0C0C080C",
		612 =>	x"08030408",
		613 =>	x"08080808",
		614 =>	x"08080403",
		615 =>	x"0C0C080C",
		616 =>	x"08030804",
		617 =>	x"04040404",
		618 =>	x"04040404",
		619 =>	x"030C080C",
		620 =>	x"08030304",
		621 =>	x"040C0C0C",
		622 =>	x"0C0C0C04",
		623 =>	x"030C080C",
		624 =>	x"08030C03",
		625 =>	x"0304040C",
		626 =>	x"04040404",
		627 =>	x"0403080C",
		628 =>	x"08030C0C",
		629 =>	x"0C030403",
		630 =>	x"0304080C",
		631 =>	x"0403080C",
		632 =>	x"08030C0C",
		633 =>	x"0C0C0304",
		634 =>	x"0404080C",
		635 =>	x"0403080C",
		636 =>	x"08030C0C",
		637 =>	x"0C0C0C03",
		638 =>	x"03040C0C",
		639 =>	x"0403080C",
		640 =>	x"08030C0C",
		641 =>	x"0C0C0C0C",
		642 =>	x"0C040404",
		643 =>	x"0403080C",
		644 =>	x"08030C0C",
		645 =>	x"0C0C0C0C",
		646 =>	x"0C030303",
		647 =>	x"030C080C",
		648 =>	x"04080808",
		649 =>	x"08080808",
		650 =>	x"08080808",
		651 =>	x"0808040C",
		652 =>	x"030C0C0C",
		653 =>	x"0C0C0C0C",
		654 =>	x"0C0C0C0C",
		655 =>	x"0C0C0C03",
		656 =>	x"03030303", -- IMG_16x16_BONUS_SHELL
		657 =>	x"03030303",
		658 =>	x"03030303",
		659 =>	x"03030303",
		660 =>	x"03080808",
		661 =>	x"08080808",
		662 =>	x"08080808",
		663 =>	x"08080403",
		664 =>	x"08030303",
		665 =>	x"03030303",
		666 =>	x"03030303",
		667 =>	x"0303080C",
		668 =>	x"08030C0C",
		669 =>	x"0C0C0C0C",
		670 =>	x"0C0C0C0C",
		671 =>	x"0C0C080C",
		672 =>	x"08030C0C",
		673 =>	x"0C0C0C0C",
		674 =>	x"0C0C0C0C",
		675 =>	x"0C0C080C",
		676 =>	x"08030C0C",
		677 =>	x"0C080808",
		678 =>	x"0404030C",
		679 =>	x"0C0C080C",
		680 =>	x"08030C0C",
		681 =>	x"08080404",
		682 =>	x"04040403",
		683 =>	x"0C0C080C",
		684 =>	x"08030C0C",
		685 =>	x"08040404",
		686 =>	x"04040403",
		687 =>	x"0C0C080C",
		688 =>	x"08030C0C",
		689 =>	x"04040404",
		690 =>	x"04040403",
		691 =>	x"0C0C080C",
		692 =>	x"08030C04",
		693 =>	x"04040404",
		694 =>	x"04040403",
		695 =>	x"0C0C080C",
		696 =>	x"08030C03",
		697 =>	x"03030303",
		698 =>	x"04040404",
		699 =>	x"030C080C",
		700 =>	x"08030C0C",
		701 =>	x"0C0C0C0C",
		702 =>	x"03030303",
		703 =>	x"030C080C",
		704 =>	x"08030C0C",
		705 =>	x"0C0C0C0C",
		706 =>	x"0C0C0C0C",
		707 =>	x"0C0C080C",
		708 =>	x"08030C0C",
		709 =>	x"0C0C0C0C",
		710 =>	x"0C0C0C0C",
		711 =>	x"0C0C080C",
		712 =>	x"04080808",
		713 =>	x"08080808",
		714 =>	x"08080808",
		715 =>	x"0808040C",
		716 =>	x"030C0C0C",
		717 =>	x"0C0C0C0C",
		718 =>	x"0C0C0C0C",
		719 =>	x"0C0C0C03",
		720 =>	x"03030303", -- IMG_16x16_BONUS_SHOVEL
		721 =>	x"03030303",
		722 =>	x"03030303",
		723 =>	x"03030303",
		724 =>	x"03080808",
		725 =>	x"08080808",
		726 =>	x"08080808",
		727 =>	x"08080403",
		728 =>	x"08030303",
		729 =>	x"03030303",
		730 =>	x"03030303",
		731 =>	x"0303080C",
		732 =>	x"08030C0C",
		733 =>	x"0C0C0C0C",
		734 =>	x"0C0C080C",
		735 =>	x"0C0C080C",
		736 =>	x"08030C0C",
		737 =>	x"0C0C0C0C",
		738 =>	x"0C0C0804",
		739 =>	x"0C0C080C",
		740 =>	x"08030C0C",
		741 =>	x"0C0C0C0C",
		742 =>	x"0C0C0404",
		743 =>	x"040C080C",
		744 =>	x"08030C0C",
		745 =>	x"0C0C0C0C",
		746 =>	x"0C080303",
		747 =>	x"030C080C",
		748 =>	x"08030C0C",
		749 =>	x"0C080C0C",
		750 =>	x"08030C0C",
		751 =>	x"0C0C080C",
		752 =>	x"08030C0C",
		753 =>	x"08080408",
		754 =>	x"030C0C0C",
		755 =>	x"0C0C080C",
		756 =>	x"08030C08",
		757 =>	x"08040C04",
		758 =>	x"030C0C0C",
		759 =>	x"0C0C080C",
		760 =>	x"08030C08",
		761 =>	x"040C0404",
		762 =>	x"04030C0C",
		763 =>	x"0C0C080C",
		764 =>	x"08030C04",
		765 =>	x"04040404",
		766 =>	x"030C0C0C",
		767 =>	x"0C0C080C",
		768 =>	x"08030C04",
		769 =>	x"04040403",
		770 =>	x"0C0C0C0C",
		771 =>	x"0C0C080C",
		772 =>	x"08030C03",
		773 =>	x"0303030C",
		774 =>	x"0C0C0C0C",
		775 =>	x"0C0C080C",
		776 =>	x"04080808",
		777 =>	x"08080808",
		778 =>	x"08080808",
		779 =>	x"0808040C",
		780 =>	x"030C0C0C",
		781 =>	x"0C0C0C0C",
		782 =>	x"0C0C0C0C",
		783 =>	x"0C0C0C03",
		784 =>	x"03030303", -- IMG_16x16_BONUS_STAR
		785 =>	x"03030303",
		786 =>	x"03030303",
		787 =>	x"03030303",
		788 =>	x"03080808",
		789 =>	x"08080808",
		790 =>	x"08080808",
		791 =>	x"08080403",
		792 =>	x"08030303",
		793 =>	x"03030303",
		794 =>	x"03030303",
		795 =>	x"0303080C",
		796 =>	x"08030C0C",
		797 =>	x"0C0C0C08",
		798 =>	x"030C0C0C",
		799 =>	x"0C0C080C",
		800 =>	x"08030C0C",
		801 =>	x"0C0C0808",
		802 =>	x"04030C0C",
		803 =>	x"0C0C080C",
		804 =>	x"08030C0C",
		805 =>	x"0C0C0808",
		806 =>	x"04030C0C",
		807 =>	x"0C0C080C",
		808 =>	x"08030808",
		809 =>	x"08080804",
		810 =>	x"04080808",
		811 =>	x"0803080C",
		812 =>	x"08030C04",
		813 =>	x"04040804",
		814 =>	x"08040404",
		815 =>	x"0303080C",
		816 =>	x"08030C0C",
		817 =>	x"04080808",
		818 =>	x"08040403",
		819 =>	x"030C080C",
		820 =>	x"08030C0C",
		821 =>	x"08080404",
		822 =>	x"08080403",
		823 =>	x"0C0C080C",
		824 =>	x"08030C04",
		825 =>	x"08040403",
		826 =>	x"04040804",
		827 =>	x"030C080C",
		828 =>	x"08030C08",
		829 =>	x"04040303",
		830 =>	x"03040408",
		831 =>	x"030C080C",
		832 =>	x"08030C04",
		833 =>	x"0303030C",
		834 =>	x"0C030304",
		835 =>	x"030C080C",
		836 =>	x"08030C03",
		837 =>	x"030C0C0C",
		838 =>	x"0C0C0C03",
		839 =>	x"030C080C",
		840 =>	x"04080808",
		841 =>	x"08080808",
		842 =>	x"08080808",
		843 =>	x"0808040C",
		844 =>	x"030C0C0C",
		845 =>	x"0C0C0C0C",
		846 =>	x"0C0C0C0C",
		847 =>	x"0C0C0C03",
		848 =>	x"03030303", -- IMG_16x16_BONUS_TANK
		849 =>	x"03030303",
		850 =>	x"03030303",
		851 =>	x"03030303",
		852 =>	x"03080808",
		853 =>	x"08080808",
		854 =>	x"08080808",
		855 =>	x"08080403",
		856 =>	x"08030303",
		857 =>	x"03030303",
		858 =>	x"03030303",
		859 =>	x"0303080C",
		860 =>	x"08030C0C",
		861 =>	x"0C0C0C0C",
		862 =>	x"0C0C0C0C",
		863 =>	x"0C0C080C",
		864 =>	x"08030C08",
		865 =>	x"0C0C0C0C",
		866 =>	x"0C0C0C0C",
		867 =>	x"0C0C080C",
		868 =>	x"08030408",
		869 =>	x"08080808",
		870 =>	x"08080403",
		871 =>	x"0C0C080C",
		872 =>	x"08030804",
		873 =>	x"04040404",
		874 =>	x"04040404",
		875 =>	x"030C080C",
		876 =>	x"08030304",
		877 =>	x"040C0C0C",
		878 =>	x"0C0C0C04",
		879 =>	x"030C080C",
		880 =>	x"08030C03",
		881 =>	x"0304040C",
		882 =>	x"04040404",
		883 =>	x"0403080C",
		884 =>	x"08030C0C",
		885 =>	x"0C030403",
		886 =>	x"0304080C",
		887 =>	x"0403080C",
		888 =>	x"08030C0C",
		889 =>	x"0C0C0304",
		890 =>	x"0404080C",
		891 =>	x"0403080C",
		892 =>	x"08030C0C",
		893 =>	x"0C0C0C03",
		894 =>	x"03040C0C",
		895 =>	x"0403080C",
		896 =>	x"08030C0C",
		897 =>	x"0C0C0C0C",
		898 =>	x"0C040404",
		899 =>	x"0403080C",
		900 =>	x"08030C0C",
		901 =>	x"0C0C0C0C",
		902 =>	x"0C030303",
		903 =>	x"030C080C",
		904 =>	x"04080808",
		905 =>	x"08080808",
		906 =>	x"08080808",
		907 =>	x"0808040C",
		908 =>	x"030C0C0C",
		909 =>	x"0C0C0C0C",
		910 =>	x"0C0C0C0C",
		911 =>	x"0C0C0C03",
		912 =>	x"03030303", -- IMG_16x16_BONUS_TIME
		913 =>	x"03030303",
		914 =>	x"03030303",
		915 =>	x"03030303",
		916 =>	x"03030808",
		917 =>	x"08080808",
		918 =>	x"08080808",
		919 =>	x"08080804",
		920 =>	x"0C080303",
		921 =>	x"03030303",
		922 =>	x"03030303",
		923 =>	x"03030308",
		924 =>	x"0C08030C",
		925 =>	x"0C0C0C08",
		926 =>	x"04080403",
		927 =>	x"0C0C0C08",
		928 =>	x"0C08030C",
		929 =>	x"0C0C0C04",
		930 =>	x"03030308",
		931 =>	x"04030C08",
		932 =>	x"0C08030C",
		933 =>	x"0C0C0404",
		934 =>	x"04040303",
		935 =>	x"03030C08",
		936 =>	x"0C08030C",
		937 =>	x"0C040808",
		938 =>	x"08080403",
		939 =>	x"0C0C0C08",
		940 =>	x"0C08030C",
		941 =>	x"0408080C",
		942 =>	x"08080804",
		943 =>	x"030C0C08",
		944 =>	x"0C08030C",
		945 =>	x"0408080C",
		946 =>	x"08080804",
		947 =>	x"030C0C08",
		948 =>	x"0C08030C",
		949 =>	x"04080808",
		950 =>	x"0C080804",
		951 =>	x"030C0C08",
		952 =>	x"0C08030C",
		953 =>	x"03040808",
		954 =>	x"08080403",
		955 =>	x"0C0C0C08",
		956 =>	x"0C08030C",
		957 =>	x"0C030404",
		958 =>	x"0404030C",
		959 =>	x"0C0C0C08",
		960 =>	x"0C08030C",
		961 =>	x"0C0C0303",
		962 =>	x"03030C0C",
		963 =>	x"0C0C0C08",
		964 =>	x"0C08030C",
		965 =>	x"0C0C0C0C",
		966 =>	x"0C0C0C0C",
		967 =>	x"0C0C0C08",
		968 =>	x"0C040808",
		969 =>	x"08080808",
		970 =>	x"08080808",
		971 =>	x"08080804",
		972 =>	x"03030C0C",
		973 =>	x"0C0C0C0C",
		974 =>	x"0C0C0C0C",
		975 =>	x"0C0C0C0C",
		976 =>	x"03030303", -- IMG_16x16_ENEMY_TANK1
		977 =>	x"03030303",
		978 =>	x"03030303",
		979 =>	x"03030303",
		980 =>	x"03030303",
		981 =>	x"03030308",
		982 =>	x"03030303",
		983 =>	x"03030303",
		984 =>	x"03030303",
		985 =>	x"03030308",
		986 =>	x"03030303",
		987 =>	x"03030303",
		988 =>	x"03030303",
		989 =>	x"03030308",
		990 =>	x"03030303",
		991 =>	x"03030303",
		992 =>	x"03080404",
		993 =>	x"03030408",
		994 =>	x"0C030308",
		995 =>	x"04040303",
		996 =>	x"030C0C04",
		997 =>	x"03080408",
		998 =>	x"0C0C0304",
		999 =>	x"0C0C0303",
		1000 =>	x"03080404",
		1001 =>	x"08080408",
		1002 =>	x"0C0C0C04",
		1003 =>	x"04040303",
		1004 =>	x"030C0C04",
		1005 =>	x"08080404",
		1006 =>	x"040C0C04",
		1007 =>	x"0C0C0303",
		1008 =>	x"03080404",
		1009 =>	x"0804040C",
		1010 =>	x"04040C04",
		1011 =>	x"04040303",
		1012 =>	x"030C0C04",
		1013 =>	x"08040C0C",
		1014 =>	x"08040C04",
		1015 =>	x"0C0C0303",
		1016 =>	x"03080404",
		1017 =>	x"08040C08",
		1018 =>	x"08040C04",
		1019 =>	x"04040303",
		1020 =>	x"030C0C04",
		1021 =>	x"08040404",
		1022 =>	x"04040C04",
		1023 =>	x"0C0C0303",
		1024 =>	x"03080404",
		1025 =>	x"08080404",
		1026 =>	x"040C0C04",
		1027 =>	x"04040303",
		1028 =>	x"030C0C04",
		1029 =>	x"03080404",
		1030 =>	x"0C0C0304",
		1031 =>	x"0C0C0303",
		1032 =>	x"03080404",
		1033 =>	x"03030C0C",
		1034 =>	x"0C030304",
		1035 =>	x"04040303",
		1036 =>	x"03030303",
		1037 =>	x"03030304",
		1038 =>	x"03030303",
		1039 =>	x"03030303",
		1040 =>	x"03030303", -- IMG_16x16_ENEMY_TANK2
		1041 =>	x"03030303",
		1042 =>	x"03030303",
		1043 =>	x"03030303",
		1044 =>	x"03030303",
		1045 =>	x"03030308",
		1046 =>	x"03030303",
		1047 =>	x"03030303",
		1048 =>	x"03030303",
		1049 =>	x"03030308",
		1050 =>	x"03030303",
		1051 =>	x"03030303",
		1052 =>	x"03040C03",
		1053 =>	x"08080C08",
		1054 =>	x"0C040403",
		1055 =>	x"040C0303",
		1056 =>	x"030C0C08",
		1057 =>	x"08080C08",
		1058 =>	x"0C040404",
		1059 =>	x"0C0C0303",
		1060 =>	x"030C0C04",
		1061 =>	x"08080C08",
		1062 =>	x"0C0C0C04",
		1063 =>	x"0C0C0303",
		1064 =>	x"03030304",
		1065 =>	x"04080408",
		1066 =>	x"040C0C04",
		1067 =>	x"03030303",
		1068 =>	x"03030304",
		1069 =>	x"08040404",
		1070 =>	x"04040C04",
		1071 =>	x"03030303",
		1072 =>	x"03040C04",
		1073 =>	x"0804040C",
		1074 =>	x"04040C04",
		1075 =>	x"040C0303",
		1076 =>	x"030C0C04",
		1077 =>	x"08040C0C",
		1078 =>	x"08040C04",
		1079 =>	x"0C0C0303",
		1080 =>	x"030C0C04",
		1081 =>	x"08040C08",
		1082 =>	x"08040C04",
		1083 =>	x"0C0C0303",
		1084 =>	x"03030304",
		1085 =>	x"08040404",
		1086 =>	x"04040C04",
		1087 =>	x"03030303",
		1088 =>	x"03030304",
		1089 =>	x"08080404",
		1090 =>	x"04080C04",
		1091 =>	x"03030303",
		1092 =>	x"03040C04",
		1093 =>	x"04040808",
		1094 =>	x"080C0C04",
		1095 =>	x"040C0303",
		1096 =>	x"030C0C04",
		1097 =>	x"0C0C0C0C",
		1098 =>	x"0C0C0C04",
		1099 =>	x"0C0C0303",
		1100 =>	x"030C0C03",
		1101 =>	x"0C0C0C08",
		1102 =>	x"0C0C0C03",
		1103 =>	x"0C0C0303",
		1104 =>	x"03030303", -- IMG_16x16_ENEMY_TANK3
		1105 =>	x"03030303",
		1106 =>	x"03030303",
		1107 =>	x"03030303",
		1108 =>	x"03030303",
		1109 =>	x"03030808",
		1110 =>	x"04030303",
		1111 =>	x"03030303",
		1112 =>	x"03030303",
		1113 =>	x"03030308",
		1114 =>	x"03030303",
		1115 =>	x"03030303",
		1116 =>	x"03030303",
		1117 =>	x"03030308",
		1118 =>	x"03030303",
		1119 =>	x"03030303",
		1120 =>	x"03080404",
		1121 =>	x"03030408",
		1122 =>	x"0C030308",
		1123 =>	x"04040303",
		1124 =>	x"030C0C04",
		1125 =>	x"03080408",
		1126 =>	x"0C0C0304",
		1127 =>	x"0C0C0303",
		1128 =>	x"03080404",
		1129 =>	x"08080408",
		1130 =>	x"0C0C0C04",
		1131 =>	x"04040303",
		1132 =>	x"030C0C04",
		1133 =>	x"08080404",
		1134 =>	x"040C0C04",
		1135 =>	x"0C0C0303",
		1136 =>	x"03080404",
		1137 =>	x"0804040C",
		1138 =>	x"04040C04",
		1139 =>	x"04040303",
		1140 =>	x"030C0C04",
		1141 =>	x"08040C0C",
		1142 =>	x"08040C04",
		1143 =>	x"0C0C0303",
		1144 =>	x"03080404",
		1145 =>	x"08040C08",
		1146 =>	x"08040C04",
		1147 =>	x"04040303",
		1148 =>	x"030C0C04",
		1149 =>	x"08040404",
		1150 =>	x"04040C04",
		1151 =>	x"0C0C0303",
		1152 =>	x"03080404",
		1153 =>	x"08080404",
		1154 =>	x"040C0C04",
		1155 =>	x"04040303",
		1156 =>	x"030C0C04",
		1157 =>	x"03080804",
		1158 =>	x"0C0C0304",
		1159 =>	x"0C0C0303",
		1160 =>	x"03080404",
		1161 =>	x"0308080C",
		1162 =>	x"0C0C0304",
		1163 =>	x"04040303",
		1164 =>	x"030C0C04",
		1165 =>	x"03030408",
		1166 =>	x"0C030304",
		1167 =>	x"0C0C0303",
		1168 =>	x"03030303", -- IMG_16x16_ENEMY_TANK4
		1169 =>	x"03030303",
		1170 =>	x"03030303",
		1171 =>	x"03030303",
		1172 =>	x"03080404",
		1173 =>	x"03030808",
		1174 =>	x"04030308",
		1175 =>	x"04040303",
		1176 =>	x"030C0C04",
		1177 =>	x"040C0808",
		1178 =>	x"040C0404",
		1179 =>	x"0C0C0303",
		1180 =>	x"03080404",
		1181 =>	x"04040408",
		1182 =>	x"0C040404",
		1183 =>	x"04040303",
		1184 =>	x"030C0C04",
		1185 =>	x"08040408",
		1186 =>	x"0C04040C",
		1187 =>	x"0C0C0303",
		1188 =>	x"03080404",
		1189 =>	x"08040408",
		1190 =>	x"0C08040C",
		1191 =>	x"04040303",
		1192 =>	x"030C0C04",
		1193 =>	x"08080408",
		1194 =>	x"0C080C0C",
		1195 =>	x"0C0C0303",
		1196 =>	x"03080404",
		1197 =>	x"08080808",
		1198 =>	x"08080C0C",
		1199 =>	x"04040303",
		1200 =>	x"030C0C04",
		1201 =>	x"0804040C",
		1202 =>	x"04040C0C",
		1203 =>	x"0C0C0303",
		1204 =>	x"03080404",
		1205 =>	x"08040C0C",
		1206 =>	x"08040C0C",
		1207 =>	x"04040303",
		1208 =>	x"030C0C04",
		1209 =>	x"08040C08",
		1210 =>	x"08040C0C",
		1211 =>	x"0C0C0303",
		1212 =>	x"03080404",
		1213 =>	x"08040404",
		1214 =>	x"04040C0C",
		1215 =>	x"04040303",
		1216 =>	x"030C0C04",
		1217 =>	x"08040404",
		1218 =>	x"04040C0C",
		1219 =>	x"0C0C0303",
		1220 =>	x"03080404",
		1221 =>	x"040C0C0C",
		1222 =>	x"0C0C040C",
		1223 =>	x"04040303",
		1224 =>	x"030C0C04",
		1225 =>	x"0C0C0C0C",
		1226 =>	x"0C0C0C04",
		1227 =>	x"0C0C0303",
		1228 =>	x"03080404",
		1229 =>	x"03030304",
		1230 =>	x"0303030C",
		1231 =>	x"04040303",
		1232 =>	x"03030303", -- IMG_16x16_EXPLOSION
		1233 =>	x"0D030D03",
		1234 =>	x"0303030D",
		1235 =>	x"03030D03",
		1236 =>	x"03080303",
		1237 =>	x"03080303",
		1238 =>	x"08030D03",
		1239 =>	x"03080D03",
		1240 =>	x"030D0D08",
		1241 =>	x"08030308",
		1242 =>	x"08030303",
		1243 =>	x"080D0303",
		1244 =>	x"03030D0D",
		1245 =>	x"080D0D08",
		1246 =>	x"0D0D0308",
		1247 =>	x"080D0303",
		1248 =>	x"0303030D",
		1249 =>	x"0E080808",
		1250 =>	x"080D0808",
		1251 =>	x"0D0D030D",
		1252 =>	x"0308030D",
		1253 =>	x"08080E08",
		1254 =>	x"0308080E",
		1255 =>	x"0D030303",
		1256 =>	x"03030D08",
		1257 =>	x"080E0D0E",
		1258 =>	x"0E030E0D",
		1259 =>	x"080D0303",
		1260 =>	x"08080808",
		1261 =>	x"03080E03",
		1262 =>	x"030E0808",
		1263 =>	x"08080808",
		1264 =>	x"030D0D0D",
		1265 =>	x"08080D0E",
		1266 =>	x"030E080D",
		1267 =>	x"0D0D0303",
		1268 =>	x"0303030D",
		1269 =>	x"0D0D0308",
		1270 =>	x"0E030D0D",
		1271 =>	x"08080303",
		1272 =>	x"03080D0D",
		1273 =>	x"08080D08",
		1274 =>	x"03080E08",
		1275 =>	x"0D0D0803",
		1276 =>	x"03030808",
		1277 =>	x"080E080D",
		1278 =>	x"080D0808",
		1279 =>	x"03030303",
		1280 =>	x"030D080D",
		1281 =>	x"0D080D08",
		1282 =>	x"080D0D08",
		1283 =>	x"08030D03",
		1284 =>	x"03080D03",
		1285 =>	x"030D030D",
		1286 =>	x"080D030D",
		1287 =>	x"0D080303",
		1288 =>	x"080D0303",
		1289 =>	x"0D030303",
		1290 =>	x"08030303",
		1291 =>	x"030D0803",
		1292 =>	x"03030303",
		1293 =>	x"03030303",
		1294 =>	x"08030D03",
		1295 =>	x"03030D03",
		1296 =>	x"03030101", -- IMG_16x16_FLAG
		1297 =>	x"01010101",
		1298 =>	x"01010101",
		1299 =>	x"01010101",
		1300 =>	x"03030202",
		1301 =>	x"01010101",
		1302 =>	x"01010101",
		1303 =>	x"01010101",
		1304 =>	x"03030202",
		1305 =>	x"02020101",
		1306 =>	x"01010101",
		1307 =>	x"01010101",
		1308 =>	x"03030202",
		1309 =>	x"02020202",
		1310 =>	x"01010101",
		1311 =>	x"01010101",
		1312 =>	x"03030202",
		1313 =>	x"02020202",
		1314 =>	x"02020101",
		1315 =>	x"01010101",
		1316 =>	x"03030202",
		1317 =>	x"02020202",
		1318 =>	x"02020202",
		1319 =>	x"01010101",
		1320 =>	x"03030202",
		1321 =>	x"02020202",
		1322 =>	x"02020202",
		1323 =>	x"02020101",
		1324 =>	x"03030202",
		1325 =>	x"02020202",
		1326 =>	x"02020202",
		1327 =>	x"02020202",
		1328 =>	x"03030202",
		1329 =>	x"02020202",
		1330 =>	x"02020202",
		1331 =>	x"02020202",
		1332 =>	x"03030101",
		1333 =>	x"01010101",
		1334 =>	x"01010101",
		1335 =>	x"01010101",
		1336 =>	x"03030101",
		1337 =>	x"01010101",
		1338 =>	x"01010101",
		1339 =>	x"01010101",
		1340 =>	x"03030101",
		1341 =>	x"01010101",
		1342 =>	x"01010101",
		1343 =>	x"01010101",
		1344 =>	x"03030101",
		1345 =>	x"01010101",
		1346 =>	x"01010101",
		1347 =>	x"01010101",
		1348 =>	x"03030101",
		1349 =>	x"01010101",
		1350 =>	x"01010101",
		1351 =>	x"01010101",
		1352 =>	x"03030101",
		1353 =>	x"01010101",
		1354 =>	x"01010101",
		1355 =>	x"01010101",
		1356 =>	x"01010101",
		1357 =>	x"01010101",
		1358 =>	x"01010101",
		1359 =>	x"01010101",
		1360 =>	x"03030303", -- IMG_16x16_MAIN_TANK
		1361 =>	x"03030303",
		1362 =>	x"03030303",
		1363 =>	x"03030303",
		1364 =>	x"03030303",
		1365 =>	x"03030303",
		1366 =>	x"03030303",
		1367 =>	x"03030303",
		1368 =>	x"03030303",
		1369 =>	x"0303030F",
		1370 =>	x"03030303",
		1371 =>	x"03030303",
		1372 =>	x"03030303",
		1373 =>	x"0303030F",
		1374 =>	x"03030303",
		1375 =>	x"03030303",
		1376 =>	x"030F1010",
		1377 =>	x"0303030F",
		1378 =>	x"0303030F",
		1379 =>	x"10100303",
		1380 =>	x"0311110F",
		1381 =>	x"0303030F",
		1382 =>	x"03030311",
		1383 =>	x"11110303",
		1384 =>	x"030F100F",
		1385 =>	x"030F100F",
		1386 =>	x"11110311",
		1387 =>	x"10100303",
		1388 =>	x"0311110F",
		1389 =>	x"0F0F1010",
		1390 =>	x"10101111",
		1391 =>	x"11110303",
		1392 =>	x"030F100F",
		1393 =>	x"0F100F0F",
		1394 =>	x"10101011",
		1395 =>	x"10100303",
		1396 =>	x"0311110F",
		1397 =>	x"0F100F10",
		1398 =>	x"11101011",
		1399 =>	x"11110303",
		1400 =>	x"030F100F",
		1401 =>	x"0F100F10",
		1402 =>	x"11101011",
		1403 =>	x"10100303",
		1404 =>	x"0311110F",
		1405 =>	x"0F0F1011",
		1406 =>	x"11101011",
		1407 =>	x"11110303",
		1408 =>	x"030F100F",
		1409 =>	x"110F0F10",
		1410 =>	x"10101111",
		1411 =>	x"10100303",
		1412 =>	x"0311110F",
		1413 =>	x"03111111",
		1414 =>	x"11110311",
		1415 =>	x"11110303",
		1416 =>	x"030F1010",
		1417 =>	x"03030303",
		1418 =>	x"03030311",
		1419 =>	x"10100303",
		1420 =>	x"03030303",
		1421 =>	x"03030303",
		1422 =>	x"03030303",
		1423 =>	x"03030303",


--			***** MAP *****


		1424 =>	x"01000100", -- z: 1 rot: 0 ptr: 256
		1425 =>	x"01000110", -- z: 1 rot: 0 ptr: 272
		1426 =>	x"01000120", -- z: 1 rot: 0 ptr: 288
		1427 =>	x"01000130", -- z: 1 rot: 0 ptr: 304
		1428 =>	x"01000140", -- z: 1 rot: 0 ptr: 320
		1429 =>	x"01000150", -- z: 1 rot: 0 ptr: 336
		1430 =>	x"01000170", -- z: 1 rot: 0 ptr: 368
		1431 =>	x"01000180", -- z: 1 rot: 0 ptr: 384
		1432 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1433 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1434 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1435 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1436 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1437 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1438 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1439 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1440 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1441 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1442 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1443 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1444 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1445 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1446 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1447 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1448 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1449 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1450 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1451 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1452 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1453 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1454 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1455 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1456 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1457 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1458 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1459 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1460 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1461 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1462 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1463 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1464 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1465 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1466 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1467 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1468 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1469 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1470 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1471 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1472 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1473 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1474 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1475 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1476 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1477 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1478 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1479 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1480 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1481 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1482 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1483 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1484 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1485 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1486 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1487 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1488 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1489 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1490 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1491 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1492 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1493 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1494 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1495 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1496 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1497 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1498 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1499 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1500 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1501 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1502 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1503 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1504 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1505 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1506 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1507 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1508 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1509 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1510 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1511 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1512 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1513 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1514 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1515 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1516 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1517 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1518 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1519 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1520 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1521 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1522 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1523 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1524 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1525 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1526 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1527 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1528 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1529 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1530 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1531 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1532 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1533 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1534 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1535 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1536 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1537 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1538 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1539 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1540 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1541 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1542 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1543 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1544 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1545 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1546 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1547 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1548 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1549 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1550 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1551 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1552 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1553 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1554 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1555 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1556 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1557 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1558 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1559 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1560 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1561 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1562 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1563 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1564 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1565 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1566 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1567 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1568 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1569 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1570 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1571 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1572 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1573 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1574 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1575 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1576 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1577 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1578 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1579 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1580 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1581 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1582 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1583 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1584 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1585 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1586 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1587 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1588 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1589 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1590 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1591 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1592 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1593 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1594 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1595 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1596 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1597 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1598 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1599 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1600 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1601 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1602 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1603 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1604 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1605 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1606 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1607 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1608 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1609 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1610 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1611 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1612 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1613 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1614 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1615 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1616 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1617 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1618 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1619 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1620 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1621 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1622 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1623 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1624 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1625 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1626 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1627 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1628 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1629 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1630 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1631 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1632 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1633 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1634 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1635 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1636 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1637 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1638 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1639 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1640 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1641 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1642 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1643 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1644 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1645 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1646 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1647 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1648 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1649 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1650 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1651 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1652 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1653 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1654 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1655 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1656 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1657 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1658 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1659 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1660 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1661 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1662 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1663 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1664 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1665 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1666 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1667 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1668 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1669 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1670 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1671 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1672 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1673 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1674 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1675 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1676 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1677 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1678 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1679 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1680 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1681 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1682 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1683 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1684 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1685 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1686 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1687 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1688 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1689 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1690 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1691 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1692 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1693 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1694 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1695 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1696 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1697 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1698 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1699 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1700 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1701 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1702 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1703 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1704 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1705 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1706 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1707 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1708 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1709 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1710 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1711 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1712 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1713 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1714 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1715 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1716 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1717 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1718 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1719 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1720 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1721 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1722 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1723 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1724 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1725 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1726 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1727 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1728 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1729 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1730 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1731 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1732 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1733 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1734 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1735 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1736 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1737 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1738 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1739 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1740 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1741 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1742 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1743 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1744 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1745 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1746 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1747 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1748 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1749 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1750 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1751 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1752 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1753 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1754 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1755 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1756 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1757 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1758 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1759 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1760 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1761 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1762 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1763 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1764 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1765 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1766 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1767 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1768 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1769 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1770 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1771 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1772 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1773 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1774 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1775 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1776 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1777 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1778 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1779 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1780 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1781 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1782 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1783 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1784 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1785 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1786 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1787 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1788 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1789 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1790 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1791 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1792 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1793 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1794 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1795 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1796 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1797 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1798 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1799 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1800 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1801 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1802 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1803 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1804 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1805 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1806 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1807 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1808 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1809 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1810 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1811 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1812 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1813 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1814 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1815 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1816 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1817 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1818 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1819 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1820 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1821 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1822 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1823 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1824 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1825 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1826 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1827 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1828 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1829 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1830 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1831 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1832 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1833 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1834 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1835 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1836 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1837 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1838 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1839 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1840 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1841 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1842 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1843 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1844 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1845 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1846 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1847 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1848 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1849 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1850 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1851 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1852 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1853 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1854 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1855 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1856 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1857 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1858 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1859 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1860 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1861 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1862 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1863 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1864 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1865 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1866 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1867 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1868 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1869 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1870 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1871 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1872 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1873 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1874 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1875 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1876 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1877 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1878 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1879 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1880 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1881 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1882 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1883 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1884 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1885 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1886 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1887 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1888 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1889 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1890 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1891 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1892 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1893 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1894 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1895 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1896 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1897 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1898 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1899 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1900 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1901 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1902 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1903 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1904 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1905 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1906 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1907 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1908 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1909 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1910 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1911 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1912 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1913 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1914 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1915 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1916 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1917 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1918 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1919 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1920 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1921 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1922 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1923 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1924 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1925 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1926 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1927 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1928 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1929 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1930 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1931 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1932 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1933 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1934 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1935 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1936 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1937 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1938 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1939 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1940 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1941 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1942 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1943 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1944 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1945 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1946 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1947 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1948 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1949 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1950 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1951 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1952 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1953 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1954 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1955 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1956 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1957 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1958 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1959 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1960 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1961 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1962 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1963 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1964 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1965 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1966 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1967 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1968 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1969 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1970 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1971 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1972 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1973 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1974 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1975 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1976 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1977 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1978 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1979 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1980 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1981 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1982 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1983 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1984 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1985 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1986 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1987 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1988 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1989 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1990 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1991 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1992 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1993 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1994 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1995 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1996 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1997 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1998 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		1999 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2000 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2001 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2002 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2003 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2004 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2005 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2006 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2007 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2008 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2009 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2010 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2011 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2012 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2013 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2014 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2015 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2016 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2017 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2018 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2019 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2020 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2021 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2022 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2023 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2024 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2025 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2026 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2027 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2028 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2029 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2030 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2031 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2032 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2033 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2034 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2035 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2036 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2037 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2038 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2039 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2040 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2041 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2042 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2043 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2044 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2045 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2046 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2047 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2048 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2049 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2050 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2051 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2052 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2053 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2054 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2055 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2056 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2057 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2058 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2059 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2060 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2061 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2062 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2063 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2064 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2065 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2066 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2067 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2068 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2069 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2070 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2071 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2072 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2073 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2074 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2075 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2076 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2077 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2078 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2079 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2080 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2081 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2082 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2083 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2084 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2085 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2086 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2087 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2088 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2089 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2090 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2091 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2092 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2093 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2094 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2095 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2096 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2097 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2098 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2099 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2100 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2101 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2102 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2103 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2104 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2105 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2106 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2107 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2108 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2109 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2110 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2111 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2112 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2113 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2114 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2115 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2116 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2117 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2118 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2119 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2120 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2121 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2122 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2123 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2124 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2125 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2126 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2127 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2128 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2129 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2130 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2131 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2132 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2133 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2134 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2135 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2136 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2137 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2138 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2139 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2140 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2141 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2142 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2143 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2144 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2145 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2146 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2147 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2148 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2149 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2150 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2151 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2152 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2153 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2154 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2155 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2156 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2157 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2158 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2159 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2160 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2161 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2162 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2163 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2164 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2165 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2166 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2167 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2168 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2169 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2170 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2171 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2172 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2173 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2174 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2175 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2176 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2177 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2178 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2179 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2180 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2181 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2182 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2183 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2184 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2185 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2186 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2187 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2188 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2189 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2190 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2191 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2192 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2193 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2194 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2195 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2196 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2197 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2198 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2199 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2200 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2201 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2202 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2203 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2204 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2205 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2206 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2207 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2208 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2209 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2210 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2211 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2212 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2213 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2214 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2215 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2216 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2217 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2218 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2219 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2220 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2221 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2222 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2223 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2224 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2225 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2226 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2227 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2228 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2229 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2230 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2231 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2232 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2233 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2234 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2235 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2236 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2237 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2238 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2239 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2240 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2241 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2242 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2243 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2244 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2245 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2246 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2247 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2248 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2249 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2250 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2251 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2252 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2253 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2254 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2255 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2256 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2257 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2258 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2259 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2260 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2261 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2262 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2263 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2264 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2265 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2266 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2267 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2268 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2269 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2270 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2271 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2272 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2273 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2274 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2275 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2276 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2277 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2278 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2279 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2280 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2281 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2282 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2283 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2284 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2285 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2286 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2287 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2288 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2289 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2290 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2291 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2292 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2293 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2294 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2295 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2296 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2297 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2298 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2299 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2300 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2301 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2302 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2303 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2304 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2305 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2306 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2307 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2308 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2309 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2310 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2311 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2312 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2313 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2314 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2315 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2316 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2317 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2318 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2319 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2320 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2321 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2322 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2323 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2324 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2325 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2326 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2327 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2328 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2329 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2330 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2331 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2332 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2333 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2334 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2335 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2336 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2337 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2338 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2339 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2340 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2341 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2342 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2343 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2344 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2345 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2346 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2347 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2348 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2349 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2350 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2351 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2352 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2353 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2354 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2355 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2356 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2357 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2358 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2359 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2360 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2361 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2362 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2363 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2364 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2365 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2366 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2367 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2368 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2369 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2370 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2371 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2372 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2373 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2374 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2375 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2376 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2377 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2378 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2379 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2380 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2381 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2382 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2383 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2384 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2385 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2386 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2387 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2388 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2389 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2390 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2391 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2392 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2393 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2394 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2395 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2396 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2397 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2398 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2399 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2400 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2401 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2402 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2403 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2404 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2405 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2406 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2407 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2408 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2409 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2410 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2411 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2412 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2413 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2414 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2415 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2416 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2417 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2418 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2419 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2420 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2421 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2422 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2423 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2424 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2425 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2426 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2427 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2428 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2429 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2430 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2431 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2432 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2433 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2434 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2435 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2436 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2437 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2438 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2439 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2440 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2441 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2442 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2443 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2444 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2445 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2446 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2447 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2448 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2449 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2450 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2451 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2452 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2453 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2454 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2455 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2456 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2457 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2458 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2459 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2460 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2461 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2462 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2463 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2464 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2465 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2466 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2467 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2468 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2469 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2470 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2471 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2472 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2473 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2474 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2475 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2476 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2477 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2478 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2479 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2480 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2481 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2482 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2483 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2484 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2485 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2486 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2487 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2488 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2489 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2490 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2491 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2492 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2493 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2494 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2495 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2496 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2497 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2498 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2499 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2500 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2501 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2502 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2503 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2504 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2505 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2506 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2507 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2508 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2509 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2510 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2511 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2512 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2513 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2514 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2515 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2516 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2517 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2518 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2519 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2520 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2521 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2522 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2523 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2524 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2525 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2526 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2527 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2528 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2529 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2530 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2531 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2532 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2533 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2534 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2535 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2536 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2537 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2538 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2539 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2540 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2541 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2542 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2543 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2544 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2545 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2546 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2547 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2548 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2549 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2550 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2551 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2552 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2553 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2554 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2555 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2556 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2557 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2558 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2559 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2560 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2561 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2562 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2563 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2564 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2565 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2566 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2567 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2568 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2569 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2570 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2571 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2572 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2573 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2574 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2575 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2576 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2577 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2578 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2579 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2580 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2581 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2582 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2583 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2584 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2585 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2586 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2587 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2588 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2589 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2590 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2591 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2592 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2593 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2594 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2595 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2596 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2597 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2598 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2599 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2600 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2601 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2602 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2603 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2604 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2605 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2606 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2607 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2608 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2609 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2610 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2611 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2612 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2613 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2614 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2615 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2616 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2617 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2618 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2619 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2620 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2621 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2622 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2623 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2624 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2625 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2626 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2627 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2628 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2629 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2630 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2631 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2632 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2633 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2634 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2635 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2636 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2637 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2638 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2639 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2640 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2641 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2642 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2643 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2644 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2645 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2646 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2647 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2648 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2649 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2650 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2651 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2652 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2653 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2654 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2655 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2656 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2657 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2658 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2659 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2660 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2661 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2662 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2663 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2664 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2665 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2666 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2667 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2668 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2669 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2670 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2671 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2672 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2673 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2674 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2675 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2676 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2677 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2678 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2679 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2680 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2681 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2682 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2683 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2684 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2685 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2686 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2687 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2688 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2689 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2690 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2691 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2692 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2693 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2694 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2695 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2696 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2697 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2698 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2699 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2700 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2701 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2702 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2703 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2704 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2705 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2706 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2707 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2708 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2709 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2710 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2711 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2712 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2713 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2714 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2715 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2716 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2717 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2718 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2719 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2720 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2721 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2722 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2723 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2724 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2725 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2726 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2727 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2728 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2729 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2730 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2731 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2732 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2733 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2734 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2735 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2736 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2737 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2738 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2739 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2740 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2741 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2742 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2743 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2744 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2745 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2746 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2747 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2748 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2749 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2750 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2751 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2752 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2753 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2754 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2755 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2756 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2757 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2758 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2759 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2760 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2761 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2762 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2763 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2764 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2765 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2766 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2767 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2768 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2769 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2770 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2771 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2772 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2773 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2774 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2775 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2776 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2777 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2778 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2779 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2780 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2781 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2782 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2783 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2784 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2785 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2786 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2787 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2788 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2789 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2790 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2791 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2792 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2793 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2794 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2795 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2796 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2797 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2798 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2799 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2800 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2801 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2802 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2803 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2804 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2805 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2806 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2807 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2808 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2809 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2810 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2811 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2812 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2813 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2814 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2815 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2816 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2817 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2818 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2819 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2820 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2821 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2822 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2823 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2824 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2825 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2826 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2827 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2828 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2829 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2830 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2831 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2832 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2833 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2834 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2835 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2836 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2837 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2838 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2839 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2840 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2841 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2842 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2843 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2844 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2845 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2846 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2847 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2848 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2849 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2850 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2851 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2852 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2853 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2854 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2855 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2856 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2857 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2858 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2859 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2860 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2861 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2862 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2863 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2864 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2865 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2866 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2867 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2868 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2869 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2870 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2871 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2872 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2873 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2874 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2875 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2876 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2877 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2878 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2879 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2880 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2881 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2882 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2883 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2884 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2885 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2886 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2887 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2888 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2889 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2890 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2891 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2892 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2893 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2894 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2895 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2896 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2897 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2898 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2899 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2900 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2901 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2902 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2903 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2904 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2905 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2906 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2907 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2908 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2909 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2910 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2911 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2912 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2913 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2914 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2915 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2916 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2917 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2918 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2919 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2920 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2921 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2922 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2923 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2924 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2925 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2926 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2927 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2928 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2929 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2930 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2931 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2932 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2933 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2934 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2935 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2936 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2937 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2938 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2939 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2940 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2941 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2942 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2943 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2944 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2945 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2946 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2947 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2948 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2949 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2950 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2951 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2952 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2953 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2954 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2955 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2956 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2957 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2958 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2959 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2960 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2961 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2962 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2963 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2964 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2965 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2966 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2967 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2968 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2969 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2970 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2971 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2972 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2973 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2974 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2975 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2976 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2977 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2978 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2979 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2980 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2981 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2982 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2983 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2984 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2985 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2986 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2987 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2988 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2989 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2990 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2991 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2992 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2993 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2994 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2995 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2996 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2997 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2998 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		2999 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3000 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3001 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3002 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3003 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3004 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3005 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3006 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3007 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3008 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3009 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3010 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3011 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3012 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3013 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3014 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3015 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3016 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3017 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3018 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3019 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3020 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3021 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3022 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3023 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3024 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3025 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3026 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3027 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3028 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3029 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3030 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3031 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3032 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3033 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3034 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3035 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3036 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3037 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3038 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3039 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3040 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3041 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3042 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3043 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3044 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3045 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3046 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3047 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3048 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3049 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3050 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3051 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3052 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3053 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3054 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3055 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3056 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3057 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3058 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3059 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3060 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3061 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3062 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3063 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3064 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3065 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3066 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3067 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3068 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3069 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3070 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3071 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3072 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3073 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3074 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3075 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3076 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3077 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3078 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3079 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3080 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3081 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3082 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3083 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3084 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3085 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3086 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3087 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3088 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3089 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3090 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3091 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3092 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3093 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3094 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3095 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3096 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3097 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3098 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3099 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3100 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3101 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3102 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3103 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3104 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3105 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3106 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3107 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3108 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3109 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3110 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3111 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3112 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3113 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3114 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3115 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3116 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3117 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3118 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3119 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3120 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3121 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3122 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3123 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3124 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3125 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3126 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3127 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3128 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3129 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3130 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3131 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3132 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3133 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3134 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3135 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3136 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3137 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3138 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3139 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3140 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3141 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3142 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3143 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3144 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3145 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3146 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3147 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3148 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3149 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3150 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3151 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3152 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3153 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3154 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3155 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3156 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3157 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3158 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3159 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3160 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3161 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3162 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3163 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3164 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3165 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3166 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3167 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3168 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3169 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3170 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3171 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3172 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3173 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3174 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3175 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3176 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3177 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3178 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3179 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3180 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3181 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3182 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3183 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3184 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3185 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3186 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3187 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3188 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3189 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3190 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3191 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3192 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3193 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3194 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3195 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3196 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3197 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3198 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3199 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3200 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3201 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3202 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3203 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3204 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3205 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3206 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3207 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3208 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3209 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3210 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3211 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3212 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3213 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3214 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3215 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3216 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3217 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3218 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3219 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3220 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3221 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3222 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3223 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3224 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3225 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3226 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3227 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3228 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3229 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3230 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3231 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3232 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3233 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3234 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3235 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3236 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3237 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3238 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3239 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3240 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3241 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3242 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3243 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3244 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3245 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3246 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3247 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3248 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3249 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3250 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3251 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3252 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3253 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3254 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3255 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3256 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3257 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3258 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3259 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3260 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3261 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3262 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3263 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3264 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3265 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3266 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3267 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3268 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3269 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3270 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3271 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3272 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3273 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3274 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3275 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3276 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3277 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3278 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3279 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3280 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3281 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3282 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3283 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3284 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3285 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3286 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3287 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3288 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3289 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3290 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3291 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3292 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3293 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3294 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3295 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3296 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3297 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3298 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3299 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3300 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3301 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3302 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3303 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3304 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3305 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3306 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3307 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3308 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3309 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3310 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3311 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3312 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3313 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3314 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3315 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3316 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3317 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3318 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3319 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3320 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3321 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3322 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3323 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3324 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3325 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3326 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3327 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3328 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3329 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3330 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3331 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3332 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3333 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3334 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3335 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3336 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3337 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3338 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3339 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3340 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3341 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3342 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3343 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3344 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3345 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3346 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3347 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3348 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3349 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3350 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3351 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3352 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3353 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3354 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3355 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3356 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3357 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3358 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3359 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3360 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3361 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3362 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3363 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3364 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3365 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3366 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3367 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3368 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3369 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3370 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3371 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3372 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3373 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3374 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3375 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3376 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3377 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3378 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3379 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3380 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3381 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3382 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3383 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3384 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3385 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3386 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3387 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3388 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3389 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3390 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3391 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3392 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3393 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3394 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3395 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3396 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3397 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3398 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3399 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3400 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3401 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3402 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3403 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3404 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3405 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3406 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3407 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3408 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3409 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3410 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3411 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3412 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3413 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3414 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3415 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3416 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3417 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3418 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3419 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3420 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3421 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3422 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3423 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3424 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3425 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3426 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3427 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3428 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3429 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3430 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3431 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3432 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3433 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3434 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3435 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3436 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3437 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3438 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3439 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3440 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3441 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3442 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3443 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3444 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3445 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3446 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3447 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3448 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3449 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3450 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3451 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3452 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3453 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3454 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3455 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3456 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3457 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3458 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3459 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3460 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3461 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3462 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3463 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3464 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3465 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3466 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3467 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3468 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3469 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3470 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3471 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3472 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3473 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3474 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3475 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3476 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3477 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3478 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3479 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3480 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3481 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3482 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3483 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3484 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3485 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3486 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3487 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3488 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3489 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3490 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3491 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3492 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3493 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3494 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3495 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3496 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3497 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3498 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3499 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3500 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3501 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3502 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3503 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3504 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3505 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3506 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3507 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3508 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3509 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3510 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3511 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3512 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3513 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3514 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3515 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3516 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3517 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3518 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3519 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3520 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3521 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3522 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3523 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3524 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3525 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3526 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3527 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3528 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3529 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3530 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3531 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3532 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3533 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3534 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3535 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3536 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3537 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3538 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3539 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3540 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3541 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3542 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3543 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3544 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3545 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3546 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3547 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3548 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3549 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3550 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3551 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3552 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3553 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3554 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3555 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3556 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3557 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3558 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3559 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3560 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3561 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3562 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3563 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3564 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3565 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3566 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3567 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3568 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3569 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3570 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3571 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3572 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3573 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3574 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3575 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3576 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3577 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3578 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3579 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3580 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3581 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3582 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3583 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3584 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3585 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3586 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3587 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3588 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3589 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3590 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3591 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3592 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3593 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3594 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3595 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3596 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3597 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3598 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3599 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3600 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3601 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3602 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3603 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3604 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3605 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3606 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3607 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3608 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3609 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3610 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3611 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3612 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3613 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3614 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3615 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3616 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3617 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3618 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3619 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3620 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3621 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3622 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3623 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3624 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3625 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3626 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3627 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3628 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3629 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3630 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3631 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3632 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3633 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3634 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3635 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3636 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3637 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3638 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3639 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3640 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3641 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3642 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3643 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3644 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3645 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3646 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3647 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3648 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3649 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3650 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3651 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3652 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3653 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3654 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3655 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3656 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3657 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3658 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3659 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3660 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3661 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3662 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3663 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3664 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3665 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3666 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3667 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3668 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3669 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3670 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3671 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3672 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3673 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3674 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3675 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3676 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3677 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3678 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3679 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3680 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3681 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3682 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3683 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3684 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3685 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3686 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3687 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3688 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3689 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3690 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3691 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3692 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3693 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3694 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3695 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3696 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3697 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3698 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3699 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3700 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3701 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3702 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3703 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3704 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3705 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3706 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3707 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3708 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3709 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3710 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3711 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3712 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3713 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3714 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3715 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3716 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3717 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3718 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3719 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3720 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3721 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3722 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3723 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3724 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3725 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3726 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3727 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3728 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3729 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3730 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3731 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3732 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3733 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3734 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3735 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3736 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3737 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3738 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3739 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3740 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3741 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3742 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3743 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3744 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3745 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3746 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3747 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3748 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3749 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3750 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3751 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3752 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3753 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3754 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3755 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3756 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3757 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3758 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3759 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3760 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3761 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3762 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3763 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3764 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3765 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3766 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3767 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3768 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3769 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3770 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3771 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3772 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3773 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3774 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3775 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3776 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3777 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3778 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3779 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3780 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3781 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3782 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3783 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3784 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3785 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3786 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3787 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3788 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3789 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3790 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3791 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3792 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3793 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3794 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3795 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3796 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3797 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3798 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3799 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3800 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3801 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3802 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3803 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3804 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3805 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3806 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3807 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3808 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3809 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3810 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3811 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3812 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3813 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3814 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3815 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3816 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3817 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3818 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3819 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3820 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3821 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3822 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3823 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3824 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3825 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3826 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3827 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3828 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3829 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3830 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3831 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3832 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3833 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3834 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3835 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3836 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3837 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3838 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3839 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3840 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3841 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3842 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3843 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3844 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3845 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3846 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3847 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3848 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3849 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3850 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3851 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3852 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3853 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3854 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3855 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3856 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3857 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3858 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3859 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3860 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3861 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3862 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3863 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3864 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3865 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3866 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3867 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3868 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3869 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3870 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3871 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3872 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3873 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3874 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3875 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3876 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3877 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3878 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3879 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3880 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3881 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3882 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3883 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3884 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3885 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3886 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3887 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3888 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3889 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3890 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3891 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3892 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3893 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3894 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3895 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3896 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3897 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3898 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3899 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3900 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3901 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3902 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3903 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3904 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3905 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3906 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3907 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3908 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3909 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3910 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3911 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3912 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3913 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3914 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3915 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3916 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3917 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3918 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3919 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3920 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3921 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3922 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3923 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3924 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3925 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3926 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3927 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3928 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3929 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3930 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3931 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3932 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3933 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3934 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3935 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3936 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3937 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3938 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3939 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3940 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3941 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3942 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3943 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3944 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3945 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3946 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3947 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3948 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3949 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3950 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3951 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3952 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3953 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3954 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3955 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3956 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3957 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3958 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3959 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3960 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3961 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3962 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3963 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3964 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3965 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3966 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3967 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3968 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3969 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3970 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3971 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3972 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3973 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3974 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3975 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3976 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3977 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3978 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3979 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3980 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3981 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3982 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3983 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3984 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3985 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3986 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3987 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3988 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3989 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3990 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3991 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3992 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3993 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3994 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3995 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3996 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3997 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3998 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		3999 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4000 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4001 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4002 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4003 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4004 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4005 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4006 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4007 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4008 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4009 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4010 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4011 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4012 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4013 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4014 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4015 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4016 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4017 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4018 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4019 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4020 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4021 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4022 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4023 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4024 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4025 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4026 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4027 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4028 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4029 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4030 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4031 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4032 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4033 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4034 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4035 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4036 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4037 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4038 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4039 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4040 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4041 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4042 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4043 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4044 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4045 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4046 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4047 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4048 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4049 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4050 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4051 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4052 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4053 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4054 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4055 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4056 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4057 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4058 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4059 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4060 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4061 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4062 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4063 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4064 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4065 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4066 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4067 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4068 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4069 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4070 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4071 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4072 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4073 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4074 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4075 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4076 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4077 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4078 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4079 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4080 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4081 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4082 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4083 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4084 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4085 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4086 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4087 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4088 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4089 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4090 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4091 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4092 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4093 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4094 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4095 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4096 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4097 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4098 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4099 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4100 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4101 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4102 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4103 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4104 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4105 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4106 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4107 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4108 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4109 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4110 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4111 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4112 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4113 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4114 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4115 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4116 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4117 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4118 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4119 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4120 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4121 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4122 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4123 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4124 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4125 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4126 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4127 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4128 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4129 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4130 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4131 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4132 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4133 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4134 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4135 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4136 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4137 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4138 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4139 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4140 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4141 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4142 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4143 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4144 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4145 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4146 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4147 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4148 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4149 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4150 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4151 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4152 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4153 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4154 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4155 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4156 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4157 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4158 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4159 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4160 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4161 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4162 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4163 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4164 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4165 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4166 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4167 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4168 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4169 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4170 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4171 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4172 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4173 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4174 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4175 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4176 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4177 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4178 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4179 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4180 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4181 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4182 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4183 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4184 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4185 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4186 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4187 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4188 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4189 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4190 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4191 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4192 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4193 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4194 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4195 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4196 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4197 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4198 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4199 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4200 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4201 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4202 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4203 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4204 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4205 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4206 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4207 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4208 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4209 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4210 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4211 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4212 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4213 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4214 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4215 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4216 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4217 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4218 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4219 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4220 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4221 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4222 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4223 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4224 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4225 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4226 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4227 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4228 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4229 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4230 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4231 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4232 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4233 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4234 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4235 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4236 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4237 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4238 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4239 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4240 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4241 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4242 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4243 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4244 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4245 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4246 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4247 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4248 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4249 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4250 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4251 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4252 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4253 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4254 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4255 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4256 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4257 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4258 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4259 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4260 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4261 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4262 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4263 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4264 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4265 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4266 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4267 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4268 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4269 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4270 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4271 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4272 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4273 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4274 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4275 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4276 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4277 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4278 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4279 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4280 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4281 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4282 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4283 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4284 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4285 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4286 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4287 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4288 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4289 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4290 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4291 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4292 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4293 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4294 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4295 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4296 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4297 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4298 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4299 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4300 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4301 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4302 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4303 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4304 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4305 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4306 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4307 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4308 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4309 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4310 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4311 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4312 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4313 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4314 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4315 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4316 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4317 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4318 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4319 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4320 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4321 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4322 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4323 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4324 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4325 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4326 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4327 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4328 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4329 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4330 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4331 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4332 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4333 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4334 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4335 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4336 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4337 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4338 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4339 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4340 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4341 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4342 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4343 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4344 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4345 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4346 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4347 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4348 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4349 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4350 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4351 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4352 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4353 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4354 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4355 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4356 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4357 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4358 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4359 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4360 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4361 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4362 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4363 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4364 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4365 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4366 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4367 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4368 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4369 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4370 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4371 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4372 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4373 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4374 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4375 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4376 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4377 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4378 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4379 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4380 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4381 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4382 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4383 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4384 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4385 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4386 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4387 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4388 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4389 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4390 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4391 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4392 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4393 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4394 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4395 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4396 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4397 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4398 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4399 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4400 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4401 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4402 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4403 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4404 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4405 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4406 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4407 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4408 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4409 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4410 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4411 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4412 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4413 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4414 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4415 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4416 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4417 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4418 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4419 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4420 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4421 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4422 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4423 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4424 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4425 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4426 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4427 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4428 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4429 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4430 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4431 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4432 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4433 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4434 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4435 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4436 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4437 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4438 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4439 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4440 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4441 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4442 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4443 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4444 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4445 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4446 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4447 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4448 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4449 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4450 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4451 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4452 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4453 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4454 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4455 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4456 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4457 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4458 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4459 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4460 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4461 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4462 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4463 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4464 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4465 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4466 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4467 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4468 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4469 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4470 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4471 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4472 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4473 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4474 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4475 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4476 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4477 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4478 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4479 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4480 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4481 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4482 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4483 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4484 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4485 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4486 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4487 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4488 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4489 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4490 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4491 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4492 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4493 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4494 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4495 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4496 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4497 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4498 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4499 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4500 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4501 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4502 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4503 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4504 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4505 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4506 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4507 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4508 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4509 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4510 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4511 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4512 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4513 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4514 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4515 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4516 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4517 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4518 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4519 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4520 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4521 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4522 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4523 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4524 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4525 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4526 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4527 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4528 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4529 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4530 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4531 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4532 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4533 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4534 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4535 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4536 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4537 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4538 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4539 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4540 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4541 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4542 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4543 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4544 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4545 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4546 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4547 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4548 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4549 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4550 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4551 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4552 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4553 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4554 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4555 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4556 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4557 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4558 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4559 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4560 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4561 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4562 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4563 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4564 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4565 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4566 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4567 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4568 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4569 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4570 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4571 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4572 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4573 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4574 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4575 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4576 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4577 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4578 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4579 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4580 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4581 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4582 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4583 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4584 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4585 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4586 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4587 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4588 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4589 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4590 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4591 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4592 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4593 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4594 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4595 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4596 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4597 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4598 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4599 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4600 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4601 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4602 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4603 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4604 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4605 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4606 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4607 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4608 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4609 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4610 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4611 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4612 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4613 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4614 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4615 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4616 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4617 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4618 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4619 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4620 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4621 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4622 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4623 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4624 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4625 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4626 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4627 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4628 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4629 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4630 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4631 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4632 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4633 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4634 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4635 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4636 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4637 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4638 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4639 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4640 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4641 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4642 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4643 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4644 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4645 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4646 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4647 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4648 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4649 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4650 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4651 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4652 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4653 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4654 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4655 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4656 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4657 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4658 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4659 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4660 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4661 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4662 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4663 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4664 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4665 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4666 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4667 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4668 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4669 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4670 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4671 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4672 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4673 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4674 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4675 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4676 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4677 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4678 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4679 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4680 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4681 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4682 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4683 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4684 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4685 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4686 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4687 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4688 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4689 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4690 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4691 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4692 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4693 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4694 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4695 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4696 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4697 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4698 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4699 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4700 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4701 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4702 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4703 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4704 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4705 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4706 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4707 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4708 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4709 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4710 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4711 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4712 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4713 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4714 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4715 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4716 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4717 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4718 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4719 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4720 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4721 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4722 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4723 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4724 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4725 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4726 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4727 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4728 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4729 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4730 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4731 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4732 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4733 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4734 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4735 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4736 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4737 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4738 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4739 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4740 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4741 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4742 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4743 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4744 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4745 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4746 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4747 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4748 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4749 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4750 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4751 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4752 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4753 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4754 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4755 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4756 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4757 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4758 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4759 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4760 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4761 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4762 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4763 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4764 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4765 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4766 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4767 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4768 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4769 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4770 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4771 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4772 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4773 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4774 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4775 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4776 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4777 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4778 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4779 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4780 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4781 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4782 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4783 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4784 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4785 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4786 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4787 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4788 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4789 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4790 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4791 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4792 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4793 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4794 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4795 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4796 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4797 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4798 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4799 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4800 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4801 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4802 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4803 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4804 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4805 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4806 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4807 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4808 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4809 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4810 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4811 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4812 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4813 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4814 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4815 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4816 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4817 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4818 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4819 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4820 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4821 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4822 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4823 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4824 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4825 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4826 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4827 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4828 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4829 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4830 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4831 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4832 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4833 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4834 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4835 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4836 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4837 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4838 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4839 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4840 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4841 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4842 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4843 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4844 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4845 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4846 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4847 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4848 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4849 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4850 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4851 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4852 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4853 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4854 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4855 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4856 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4857 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4858 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4859 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4860 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4861 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4862 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4863 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4864 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4865 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4866 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4867 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4868 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4869 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4870 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4871 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4872 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4873 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4874 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4875 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4876 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4877 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4878 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4879 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4880 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4881 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4882 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4883 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4884 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4885 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4886 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4887 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4888 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4889 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4890 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4891 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4892 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4893 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4894 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4895 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4896 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4897 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4898 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4899 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4900 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4901 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4902 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4903 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4904 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4905 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4906 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4907 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4908 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4909 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4910 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4911 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4912 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4913 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4914 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4915 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4916 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4917 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4918 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4919 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4920 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4921 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4922 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4923 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4924 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4925 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4926 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4927 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4928 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4929 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4930 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4931 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4932 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4933 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4934 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4935 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4936 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4937 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4938 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4939 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4940 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4941 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4942 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4943 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4944 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4945 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4946 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4947 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4948 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4949 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4950 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4951 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4952 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4953 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4954 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4955 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4956 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4957 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4958 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4959 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4960 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4961 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4962 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4963 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4964 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4965 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4966 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4967 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4968 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4969 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4970 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4971 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4972 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4973 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4974 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4975 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4976 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4977 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4978 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4979 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4980 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4981 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4982 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4983 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4984 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4985 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4986 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4987 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4988 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4989 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4990 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4991 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4992 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4993 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4994 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4995 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4996 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4997 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4998 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		4999 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5000 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5001 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5002 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5003 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5004 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5005 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5006 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5007 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5008 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5009 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5010 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5011 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5012 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5013 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5014 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5015 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5016 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5017 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5018 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5019 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5020 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5021 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5022 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5023 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5024 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5025 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5026 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5027 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5028 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5029 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5030 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5031 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5032 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5033 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5034 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5035 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5036 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5037 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5038 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5039 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5040 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5041 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5042 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5043 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5044 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5045 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5046 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5047 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5048 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5049 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5050 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5051 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5052 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5053 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5054 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5055 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5056 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5057 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5058 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5059 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5060 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5061 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5062 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5063 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5064 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5065 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5066 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5067 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5068 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5069 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5070 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5071 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5072 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5073 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5074 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5075 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5076 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5077 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5078 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5079 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5080 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5081 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5082 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5083 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5084 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5085 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5086 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5087 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5088 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5089 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5090 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5091 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5092 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5093 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5094 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5095 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5096 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5097 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5098 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5099 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5100 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5101 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5102 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5103 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5104 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5105 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5106 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5107 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5108 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5109 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5110 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5111 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5112 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5113 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5114 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5115 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5116 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5117 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5118 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5119 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5120 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5121 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5122 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5123 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5124 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5125 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5126 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5127 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5128 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5129 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5130 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5131 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5132 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5133 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5134 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5135 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5136 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5137 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5138 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5139 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5140 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5141 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5142 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5143 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5144 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5145 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5146 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5147 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5148 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5149 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5150 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5151 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5152 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5153 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5154 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5155 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5156 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5157 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5158 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5159 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5160 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5161 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5162 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5163 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5164 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5165 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5166 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5167 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5168 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5169 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5170 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5171 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5172 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5173 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5174 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5175 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5176 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5177 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5178 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5179 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5180 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5181 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5182 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5183 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5184 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5185 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5186 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5187 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5188 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5189 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5190 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5191 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5192 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5193 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5194 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5195 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5196 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5197 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5198 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5199 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5200 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5201 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5202 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5203 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5204 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5205 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5206 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5207 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5208 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5209 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5210 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5211 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5212 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5213 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5214 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5215 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5216 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5217 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5218 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5219 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5220 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5221 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5222 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5223 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5224 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5225 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5226 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5227 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5228 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5229 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5230 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5231 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5232 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5233 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5234 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5235 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5236 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5237 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5238 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5239 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5240 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5241 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5242 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5243 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5244 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5245 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5246 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5247 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5248 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5249 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5250 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5251 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5252 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5253 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5254 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5255 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5256 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5257 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5258 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5259 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5260 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5261 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5262 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5263 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5264 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5265 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5266 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5267 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5268 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5269 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5270 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5271 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5272 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5273 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5274 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5275 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5276 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5277 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5278 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5279 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5280 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5281 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5282 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5283 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5284 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5285 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5286 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5287 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5288 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5289 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5290 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5291 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5292 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5293 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5294 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5295 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5296 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5297 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5298 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5299 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5300 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5301 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5302 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5303 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5304 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5305 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5306 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5307 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5308 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5309 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5310 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5311 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5312 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5313 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5314 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5315 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5316 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5317 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5318 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5319 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5320 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5321 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5322 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5323 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5324 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5325 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5326 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5327 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5328 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5329 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5330 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5331 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5332 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5333 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5334 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5335 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5336 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5337 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5338 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5339 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5340 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5341 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5342 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5343 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5344 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5345 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5346 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5347 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5348 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5349 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5350 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5351 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5352 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5353 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5354 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5355 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5356 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5357 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5358 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5359 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5360 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5361 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5362 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5363 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5364 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5365 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5366 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5367 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5368 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5369 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5370 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5371 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5372 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5373 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5374 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5375 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5376 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5377 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5378 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5379 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5380 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5381 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5382 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5383 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5384 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5385 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5386 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5387 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5388 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5389 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5390 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5391 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5392 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5393 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5394 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5395 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5396 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5397 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5398 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5399 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5400 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5401 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5402 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5403 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5404 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5405 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5406 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5407 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5408 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5409 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5410 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5411 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5412 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5413 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5414 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5415 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5416 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5417 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5418 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5419 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5420 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5421 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5422 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5423 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5424 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5425 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5426 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5427 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5428 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5429 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5430 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5431 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5432 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5433 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5434 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5435 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5436 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5437 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5438 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5439 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5440 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5441 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5442 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5443 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5444 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5445 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5446 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5447 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5448 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5449 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5450 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5451 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5452 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5453 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5454 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5455 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5456 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5457 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5458 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5459 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5460 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5461 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5462 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5463 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5464 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5465 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5466 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5467 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5468 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5469 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5470 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5471 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5472 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5473 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5474 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5475 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5476 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5477 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5478 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5479 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5480 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5481 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5482 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5483 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5484 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5485 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5486 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5487 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5488 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5489 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5490 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5491 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5492 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5493 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5494 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5495 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5496 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5497 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5498 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5499 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5500 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5501 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5502 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5503 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5504 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5505 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5506 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5507 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5508 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5509 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5510 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5511 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5512 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5513 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5514 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5515 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5516 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5517 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5518 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5519 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5520 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5521 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5522 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5523 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5524 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5525 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5526 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5527 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5528 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5529 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5530 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5531 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5532 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5533 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5534 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5535 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5536 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5537 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5538 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5539 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5540 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5541 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5542 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5543 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5544 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5545 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5546 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5547 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5548 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5549 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5550 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5551 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5552 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5553 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5554 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5555 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5556 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5557 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5558 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5559 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5560 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5561 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5562 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5563 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5564 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5565 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5566 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5567 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5568 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5569 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5570 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5571 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5572 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5573 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5574 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5575 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5576 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5577 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5578 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5579 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5580 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5581 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5582 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5583 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5584 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5585 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5586 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5587 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5588 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5589 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5590 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5591 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5592 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5593 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5594 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5595 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5596 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5597 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5598 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5599 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5600 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5601 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5602 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5603 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5604 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5605 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5606 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5607 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5608 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5609 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5610 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5611 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5612 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5613 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5614 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5615 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5616 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5617 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5618 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5619 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5620 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5621 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5622 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5623 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5624 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5625 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5626 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5627 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5628 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5629 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5630 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5631 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5632 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5633 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5634 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5635 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5636 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5637 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5638 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5639 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5640 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5641 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5642 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5643 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5644 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5645 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5646 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5647 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5648 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5649 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5650 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5651 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5652 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5653 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5654 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5655 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5656 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5657 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5658 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5659 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5660 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5661 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5662 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5663 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5664 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5665 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5666 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5667 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5668 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5669 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5670 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5671 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5672 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5673 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5674 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5675 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5676 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5677 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5678 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5679 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5680 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5681 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5682 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5683 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5684 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5685 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5686 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5687 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5688 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5689 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5690 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5691 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5692 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5693 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5694 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5695 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5696 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5697 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5698 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5699 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5700 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5701 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5702 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5703 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5704 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5705 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5706 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5707 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5708 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5709 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5710 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5711 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5712 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5713 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5714 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5715 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5716 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5717 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5718 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5719 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5720 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5721 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5722 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5723 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5724 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5725 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5726 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5727 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5728 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5729 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5730 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5731 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5732 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5733 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5734 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5735 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5736 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5737 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5738 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5739 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5740 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5741 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5742 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5743 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5744 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5745 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5746 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5747 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5748 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5749 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5750 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5751 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5752 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5753 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5754 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5755 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5756 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5757 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5758 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5759 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5760 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5761 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5762 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5763 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5764 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5765 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5766 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5767 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5768 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5769 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5770 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5771 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5772 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5773 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5774 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5775 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5776 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5777 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5778 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5779 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5780 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5781 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5782 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5783 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5784 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5785 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5786 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5787 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5788 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5789 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5790 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5791 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5792 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5793 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5794 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5795 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5796 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5797 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5798 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5799 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5800 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5801 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5802 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5803 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5804 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5805 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5806 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5807 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5808 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5809 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5810 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5811 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5812 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5813 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5814 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5815 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5816 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5817 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5818 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5819 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5820 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5821 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5822 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5823 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5824 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5825 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5826 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5827 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5828 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5829 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5830 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5831 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5832 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5833 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5834 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5835 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5836 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5837 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5838 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5839 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5840 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5841 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5842 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5843 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5844 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5845 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5846 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5847 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5848 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5849 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5850 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5851 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5852 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5853 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5854 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5855 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5856 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5857 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5858 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5859 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5860 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5861 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5862 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5863 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5864 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5865 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5866 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5867 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5868 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5869 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5870 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5871 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5872 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5873 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5874 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5875 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5876 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5877 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5878 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5879 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5880 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5881 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5882 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5883 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5884 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5885 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5886 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5887 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5888 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5889 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5890 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5891 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5892 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5893 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5894 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5895 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5896 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5897 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5898 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5899 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5900 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5901 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5902 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5903 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5904 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5905 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5906 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5907 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5908 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5909 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5910 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5911 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5912 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5913 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5914 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5915 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5916 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5917 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5918 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5919 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5920 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5921 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5922 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5923 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5924 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5925 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5926 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5927 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5928 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5929 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5930 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5931 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5932 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5933 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5934 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5935 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5936 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5937 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5938 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5939 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5940 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5941 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5942 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5943 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5944 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5945 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5946 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5947 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5948 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5949 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5950 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5951 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5952 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5953 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5954 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5955 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5956 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5957 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5958 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5959 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5960 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5961 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5962 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5963 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5964 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5965 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5966 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5967 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5968 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5969 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5970 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5971 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5972 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5973 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5974 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5975 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5976 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5977 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5978 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5979 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5980 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5981 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5982 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5983 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5984 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5985 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5986 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5987 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5988 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5989 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5990 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5991 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5992 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5993 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5994 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5995 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5996 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5997 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5998 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		5999 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6000 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6001 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6002 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6003 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6004 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6005 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6006 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6007 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6008 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6009 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6010 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6011 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6012 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6013 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6014 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6015 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6016 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6017 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6018 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6019 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6020 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6021 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6022 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6023 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6024 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6025 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6026 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6027 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6028 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6029 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6030 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6031 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6032 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6033 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6034 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6035 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6036 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6037 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6038 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6039 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6040 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6041 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6042 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6043 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6044 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6045 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6046 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6047 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6048 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6049 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6050 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6051 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6052 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6053 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6054 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6055 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6056 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6057 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6058 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6059 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6060 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6061 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6062 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6063 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6064 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6065 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6066 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6067 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6068 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6069 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6070 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6071 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6072 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6073 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6074 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6075 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6076 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6077 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6078 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6079 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6080 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6081 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6082 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6083 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6084 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6085 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6086 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6087 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6088 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6089 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6090 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6091 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6092 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6093 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6094 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6095 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6096 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6097 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6098 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6099 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6100 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6101 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6102 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6103 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6104 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6105 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6106 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6107 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6108 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6109 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6110 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6111 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6112 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6113 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6114 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6115 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6116 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6117 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6118 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6119 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6120 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6121 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6122 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6123 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6124 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6125 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6126 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6127 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6128 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6129 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6130 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6131 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6132 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6133 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6134 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6135 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6136 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6137 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6138 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6139 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6140 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6141 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6142 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6143 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6144 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6145 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6146 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6147 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6148 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6149 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6150 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6151 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6152 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6153 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6154 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6155 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6156 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6157 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6158 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6159 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6160 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6161 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6162 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6163 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6164 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6165 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6166 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6167 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6168 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6169 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6170 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6171 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6172 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6173 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6174 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6175 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6176 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6177 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6178 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6179 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6180 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6181 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6182 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6183 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6184 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6185 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6186 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6187 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6188 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6189 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6190 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6191 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6192 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6193 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6194 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6195 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6196 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6197 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6198 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6199 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6200 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6201 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6202 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6203 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6204 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6205 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6206 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6207 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6208 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6209 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6210 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6211 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6212 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6213 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6214 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6215 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6216 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6217 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6218 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6219 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6220 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6221 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6222 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		6223 =>	x"00000160", -- z: 0 rot: 0 ptr: 352
		others => x"00000000"
	);

begin

	process(clk_i) begin
		if rising_edge(clk_i) then
--			if we_i = '1' then
--				mem( to_integer( unsigned( addr_i ) ) ) <= data_o;
--			end if;
			data_o <= mem(to_integer(addr_i));
		end if; 
	end process;

end architecture arch;