
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

-- GENERATED BY BC_MEM_PACKER
-- DATE: Fri Jul 10 13:01:11 2015

	signal mem : ram_t := (


--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00808000", -- R: 0 G: 128 B: 128
		2 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		3 =>	x"00000080", -- R: 128 G: 0 B: 0
		4 =>	x"00806060", -- R: 96 G: 96 B: 128
		5 =>	x"000040A0", -- R: 160 G: 64 B: 0
		6 =>	x"00006000", -- R: 0 G: 96 B: 0
		7 =>	x"00004000", -- R: 0 G: 64 B: 0
		8 =>	x"0000E080", -- R: 128 G: 224 B: 0
		9 =>	x"00A4A0A0", -- R: 160 G: 160 B: 164
		10 =>	x"00C04040", -- R: 64 G: 64 B: 192
		11 =>	x"00F0CAA6", -- R: 166 G: 202 B: 240
		12 =>	x"00404000", -- R: 0 G: 64 B: 64
		13 =>	x"00800060", -- R: 96 G: 0 B: 128
		14 =>	x"004040C0", -- R: 192 G: 64 B: 64
		15 =>	x"0080E0E0", -- R: 224 G: 224 B: 128
		16 =>	x"0040A0E0", -- R: 224 G: 160 B: 64
		17 =>	x"00006060", -- R: 96 G: 96 B: 0
		18 =>	x"00000000", -- Unused
		19 =>	x"00000000", -- Unused
		20 =>	x"00000000", -- Unused
		21 =>	x"00000000", -- Unused
		22 =>	x"00000000", -- Unused
		23 =>	x"00000000", -- Unused
		24 =>	x"00000000", -- Unused
		25 =>	x"00000000", -- Unused
		26 =>	x"00000000", -- Unused
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused


--			***** 8x8 IMAGES *****


		256 =>	x"01010101", -- IMG_8x8_01_A
		257 =>	x"01010101",
		258 =>	x"01010102",
		259 =>	x"02010101",
		260 =>	x"01010201",
		261 =>	x"01020101",
		262 =>	x"01010201",
		263 =>	x"01020101",
		264 =>	x"01010202",
		265 =>	x"02020101",
		266 =>	x"01010201",
		267 =>	x"01020101",
		268 =>	x"01010201",
		269 =>	x"01020101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01010101", -- IMG_8x8_02_B
		273 =>	x"01010101",
		274 =>	x"01010202",
		275 =>	x"02020101",
		276 =>	x"01010201",
		277 =>	x"01010101",
		278 =>	x"01010202",
		279 =>	x"02010101",
		280 =>	x"01010201",
		281 =>	x"01020101",
		282 =>	x"01010201",
		283 =>	x"01020101",
		284 =>	x"01010202",
		285 =>	x"02010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01010101", -- IMG_8x8_03_V
		289 =>	x"01010101",
		290 =>	x"01010202",
		291 =>	x"02010101",
		292 =>	x"01010201",
		293 =>	x"01020101",
		294 =>	x"01010201",
		295 =>	x"01020101",
		296 =>	x"01010202",
		297 =>	x"02010101",
		298 =>	x"01010201",
		299 =>	x"01020101",
		300 =>	x"01010202",
		301 =>	x"02010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"01010101", -- IMG_8x8_04_G
		305 =>	x"01010101",
		306 =>	x"01010202",
		307 =>	x"02020101",
		308 =>	x"01010201",
		309 =>	x"01020101",
		310 =>	x"01010201",
		311 =>	x"01010101",
		312 =>	x"01010201",
		313 =>	x"01010101",
		314 =>	x"01010201",
		315 =>	x"01010101",
		316 =>	x"01010201",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101",
		320 =>	x"01010101", -- IMG_8x8_05_D
		321 =>	x"01010101",
		322 =>	x"01010101",
		323 =>	x"02020101",
		324 =>	x"01010102",
		325 =>	x"01020101",
		326 =>	x"01010102",
		327 =>	x"01020101",
		328 =>	x"01010102",
		329 =>	x"01020101",
		330 =>	x"01010202",
		331 =>	x"02020101",
		332 =>	x"01010201",
		333 =>	x"01020101",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"01010101", -- IMG_8x8_06_DJ
		337 =>	x"01010101",
		338 =>	x"01010202",
		339 =>	x"02020101",
		340 =>	x"01010102",
		341 =>	x"01010101",
		342 =>	x"01010102",
		343 =>	x"02010101",
		344 =>	x"01010102",
		345 =>	x"01020101",
		346 =>	x"01010101",
		347 =>	x"01020101",
		348 =>	x"01010202",
		349 =>	x"02010101",
		350 =>	x"01010101",
		351 =>	x"01010101",
		352 =>	x"01010101", -- IMG_8x8_07_E
		353 =>	x"01010101",
		354 =>	x"01010202",
		355 =>	x"02020101",
		356 =>	x"01010201",
		357 =>	x"01010101",
		358 =>	x"01010201",
		359 =>	x"01010101",
		360 =>	x"01010202",
		361 =>	x"02010101",
		362 =>	x"01010201",
		363 =>	x"01010101",
		364 =>	x"01010202",
		365 =>	x"02020101",
		366 =>	x"01010101",
		367 =>	x"01010101",
		368 =>	x"01010101", -- IMG_8x8_08_ZH
		369 =>	x"01010101",
		370 =>	x"01020102",
		371 =>	x"01020101",
		372 =>	x"01020102",
		373 =>	x"01020101",
		374 =>	x"01020202",
		375 =>	x"02020101",
		376 =>	x"01010102",
		377 =>	x"01010101",
		378 =>	x"01020202",
		379 =>	x"02020101",
		380 =>	x"01020102",
		381 =>	x"01020101",
		382 =>	x"01010101",
		383 =>	x"01010101",
		384 =>	x"01010101", -- IMG_8x8_09_Z
		385 =>	x"01010101",
		386 =>	x"01010202",
		387 =>	x"02020101",
		388 =>	x"01010201",
		389 =>	x"01020101",
		390 =>	x"01010101",
		391 =>	x"02010101",
		392 =>	x"01010102",
		393 =>	x"02020101",
		394 =>	x"01010101",
		395 =>	x"01020101",
		396 =>	x"01010202",
		397 =>	x"02020101",
		398 =>	x"01010101",
		399 =>	x"01010101",
		400 =>	x"01010101", -- IMG_8x8_10_I
		401 =>	x"01010101",
		402 =>	x"01010201",
		403 =>	x"01020101",
		404 =>	x"01010201",
		405 =>	x"01020101",
		406 =>	x"01010201",
		407 =>	x"02020101",
		408 =>	x"01010202",
		409 =>	x"01020101",
		410 =>	x"01010201",
		411 =>	x"01020101",
		412 =>	x"01010201",
		413 =>	x"01020101",
		414 =>	x"01010101",
		415 =>	x"01010101",
		416 =>	x"01010101", -- IMG_8x8_11_J
		417 =>	x"01010101",
		418 =>	x"01010202",
		419 =>	x"02020101",
		420 =>	x"01010101",
		421 =>	x"01020101",
		422 =>	x"01010101",
		423 =>	x"01020101",
		424 =>	x"01010201",
		425 =>	x"01020101",
		426 =>	x"01010201",
		427 =>	x"01020101",
		428 =>	x"01010102",
		429 =>	x"02010101",
		430 =>	x"01010101",
		431 =>	x"01010101",
		432 =>	x"01010101", -- IMG_8x8_12_K
		433 =>	x"01010101",
		434 =>	x"01010201",
		435 =>	x"01020101",
		436 =>	x"01010201",
		437 =>	x"01020101",
		438 =>	x"01010201",
		439 =>	x"02010101",
		440 =>	x"01010202",
		441 =>	x"01010101",
		442 =>	x"01010201",
		443 =>	x"02010101",
		444 =>	x"01010201",
		445 =>	x"01020101",
		446 =>	x"01010101",
		447 =>	x"01010101",
		448 =>	x"01010101", -- IMG_8x8_13_L
		449 =>	x"01010101",
		450 =>	x"01010102",
		451 =>	x"02020101",
		452 =>	x"01010201",
		453 =>	x"01020101",
		454 =>	x"01010201",
		455 =>	x"01020101",
		456 =>	x"01010201",
		457 =>	x"01020101",
		458 =>	x"01010201",
		459 =>	x"01020101",
		460 =>	x"01020201",
		461 =>	x"01020101",
		462 =>	x"01010101",
		463 =>	x"01010101",
		464 =>	x"01010101", -- IMG_8x8_14_LJ
		465 =>	x"01010101",
		466 =>	x"01010102",
		467 =>	x"02010101",
		468 =>	x"01010201",
		469 =>	x"02010101",
		470 =>	x"01010201",
		471 =>	x"02020101",
		472 =>	x"01010201",
		473 =>	x"02010201",
		474 =>	x"01010201",
		475 =>	x"02010201",
		476 =>	x"01020201",
		477 =>	x"02020101",
		478 =>	x"01010101",
		479 =>	x"01010101",
		480 =>	x"01010101", -- IMG_8x8_15_M
		481 =>	x"01010101",
		482 =>	x"01020101",
		483 =>	x"01020101",
		484 =>	x"01020201",
		485 =>	x"02020101",
		486 =>	x"01020102",
		487 =>	x"01020101",
		488 =>	x"01020101",
		489 =>	x"01020101",
		490 =>	x"01020101",
		491 =>	x"01020101",
		492 =>	x"01020101",
		493 =>	x"01020101",
		494 =>	x"01010101",
		495 =>	x"01010101",
		496 =>	x"01010101", -- IMG_8x8_16_N
		497 =>	x"01010101",
		498 =>	x"01010201",
		499 =>	x"01020101",
		500 =>	x"01010201",
		501 =>	x"01020101",
		502 =>	x"01010202",
		503 =>	x"02020101",
		504 =>	x"01010201",
		505 =>	x"01020101",
		506 =>	x"01010201",
		507 =>	x"01020101",
		508 =>	x"01010201",
		509 =>	x"01020101",
		510 =>	x"01010101",
		511 =>	x"01010101",
		512 =>	x"01010101", -- IMG_8x8_17_NJ
		513 =>	x"01010101",
		514 =>	x"01020101",
		515 =>	x"02010101",
		516 =>	x"01020101",
		517 =>	x"02010101",
		518 =>	x"01020202",
		519 =>	x"02020101",
		520 =>	x"01020101",
		521 =>	x"02010201",
		522 =>	x"01020101",
		523 =>	x"02010201",
		524 =>	x"01020101",
		525 =>	x"02020101",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"01010101", -- IMG_8x8_18_O
		529 =>	x"01010101",
		530 =>	x"01010102",
		531 =>	x"02010101",
		532 =>	x"01010201",
		533 =>	x"01020101",
		534 =>	x"01010201",
		535 =>	x"01020101",
		536 =>	x"01010201",
		537 =>	x"01020101",
		538 =>	x"01010201",
		539 =>	x"01020101",
		540 =>	x"01010102",
		541 =>	x"02010101",
		542 =>	x"01010101",
		543 =>	x"01010101",
		544 =>	x"01010101", -- IMG_8x8_19_P
		545 =>	x"01010101",
		546 =>	x"01010202",
		547 =>	x"02020101",
		548 =>	x"01010201",
		549 =>	x"01020101",
		550 =>	x"01010201",
		551 =>	x"01020101",
		552 =>	x"01010201",
		553 =>	x"01020101",
		554 =>	x"01010201",
		555 =>	x"01020101",
		556 =>	x"01010201",
		557 =>	x"01020101",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01010101", -- IMG_8x8_20_R
		561 =>	x"01010101",
		562 =>	x"01010202",
		563 =>	x"02010101",
		564 =>	x"01010201",
		565 =>	x"01020101",
		566 =>	x"01010201",
		567 =>	x"01020101",
		568 =>	x"01010202",
		569 =>	x"02010101",
		570 =>	x"01010201",
		571 =>	x"01010101",
		572 =>	x"01010201",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101",
		576 =>	x"01010101", -- IMG_8x8_21_S
		577 =>	x"01010101",
		578 =>	x"01010102",
		579 =>	x"02020101",
		580 =>	x"01010201",
		581 =>	x"01020101",
		582 =>	x"01010201",
		583 =>	x"01010101",
		584 =>	x"01010201",
		585 =>	x"01010101",
		586 =>	x"01010201",
		587 =>	x"01020101",
		588 =>	x"01010102",
		589 =>	x"02020101",
		590 =>	x"01010101",
		591 =>	x"01010101",
		592 =>	x"01010101", -- IMG_8x8_22_T
		593 =>	x"01010101",
		594 =>	x"01020202",
		595 =>	x"02020101",
		596 =>	x"01010102",
		597 =>	x"01010101",
		598 =>	x"01010102",
		599 =>	x"01010101",
		600 =>	x"01010102",
		601 =>	x"01010101",
		602 =>	x"01010102",
		603 =>	x"01010101",
		604 =>	x"01010102",
		605 =>	x"01010101",
		606 =>	x"01010101",
		607 =>	x"01010101",
		608 =>	x"01010101", -- IMG_8x8_23_TJ
		609 =>	x"01010101",
		610 =>	x"01020202",
		611 =>	x"02010101",
		612 =>	x"01010201",
		613 =>	x"01010101",
		614 =>	x"01010202",
		615 =>	x"02010101",
		616 =>	x"01010201",
		617 =>	x"01020101",
		618 =>	x"01010201",
		619 =>	x"01020101",
		620 =>	x"01010201",
		621 =>	x"01020101",
		622 =>	x"01010101",
		623 =>	x"01010101",
		624 =>	x"01010101", -- IMG_8x8_24_U
		625 =>	x"01010101",
		626 =>	x"01010201",
		627 =>	x"01020101",
		628 =>	x"01010201",
		629 =>	x"01020101",
		630 =>	x"01010201",
		631 =>	x"01020101",
		632 =>	x"01010102",
		633 =>	x"02020101",
		634 =>	x"01010101",
		635 =>	x"01020101",
		636 =>	x"01010202",
		637 =>	x"02010101",
		638 =>	x"01010101",
		639 =>	x"01010101",
		640 =>	x"01010101", -- IMG_8x8_25_F
		641 =>	x"01010101",
		642 =>	x"01010102",
		643 =>	x"01010101",
		644 =>	x"01020202",
		645 =>	x"02020101",
		646 =>	x"01020102",
		647 =>	x"01020101",
		648 =>	x"01020102",
		649 =>	x"01020101",
		650 =>	x"01020202",
		651 =>	x"02020101",
		652 =>	x"01010102",
		653 =>	x"01010101",
		654 =>	x"01010101",
		655 =>	x"01010101",
		656 =>	x"01010101", -- IMG_8x8_26_H
		657 =>	x"01010101",
		658 =>	x"01010201",
		659 =>	x"01020101",
		660 =>	x"01010201",
		661 =>	x"01020101",
		662 =>	x"01010201",
		663 =>	x"01020101",
		664 =>	x"01010102",
		665 =>	x"02010101",
		666 =>	x"01010201",
		667 =>	x"01020101",
		668 =>	x"01010201",
		669 =>	x"01020101",
		670 =>	x"01010101",
		671 =>	x"01010101",
		672 =>	x"01010101", -- IMG_8x8_27_C
		673 =>	x"01010101",
		674 =>	x"01010201",
		675 =>	x"02010101",
		676 =>	x"01010201",
		677 =>	x"02010101",
		678 =>	x"01010201",
		679 =>	x"02010101",
		680 =>	x"01010201",
		681 =>	x"02010101",
		682 =>	x"01010202",
		683 =>	x"02020101",
		684 =>	x"01010101",
		685 =>	x"01020101",
		686 =>	x"01010101",
		687 =>	x"01010101",
		688 =>	x"01010101", -- IMG_8x8_28_CH
		689 =>	x"01010101",
		690 =>	x"01010201",
		691 =>	x"01020101",
		692 =>	x"01010201",
		693 =>	x"01020101",
		694 =>	x"01010201",
		695 =>	x"01020101",
		696 =>	x"01010102",
		697 =>	x"02020101",
		698 =>	x"01010101",
		699 =>	x"01020101",
		700 =>	x"01010101",
		701 =>	x"01020101",
		702 =>	x"01010101",
		703 =>	x"01010101",
		704 =>	x"01010101", -- IMG_8x8_29_DZH
		705 =>	x"01010101",
		706 =>	x"01020101",
		707 =>	x"01020101",
		708 =>	x"01020101",
		709 =>	x"01020101",
		710 =>	x"01020101",
		711 =>	x"01020101",
		712 =>	x"01020101",
		713 =>	x"01020101",
		714 =>	x"01020202",
		715 =>	x"02020101",
		716 =>	x"01010102",
		717 =>	x"01010101",
		718 =>	x"01010101",
		719 =>	x"01010101",
		720 =>	x"01010101", -- IMG_8x8_30_SH
		721 =>	x"01010101",
		722 =>	x"01020102",
		723 =>	x"01020101",
		724 =>	x"01020102",
		725 =>	x"01020101",
		726 =>	x"01020102",
		727 =>	x"01020101",
		728 =>	x"01020102",
		729 =>	x"01020101",
		730 =>	x"01020102",
		731 =>	x"01020101",
		732 =>	x"01020202",
		733 =>	x"02020101",
		734 =>	x"01010101",
		735 =>	x"01010101",
		736 =>	x"01010101", -- IMG_8x8_31_NUM_0
		737 =>	x"01010101",
		738 =>	x"01010102",
		739 =>	x"02010101",
		740 =>	x"01010201",
		741 =>	x"01020101",
		742 =>	x"01010201",
		743 =>	x"02020101",
		744 =>	x"01010202",
		745 =>	x"01020101",
		746 =>	x"01010201",
		747 =>	x"01020101",
		748 =>	x"01010102",
		749 =>	x"02010101",
		750 =>	x"01010101",
		751 =>	x"01010101",
		752 =>	x"01010101", -- IMG_8x8_32_NUM_1
		753 =>	x"01010101",
		754 =>	x"01010102",
		755 =>	x"01010101",
		756 =>	x"01010202",
		757 =>	x"01010101",
		758 =>	x"01010102",
		759 =>	x"01010101",
		760 =>	x"01010102",
		761 =>	x"01010101",
		762 =>	x"01010102",
		763 =>	x"01010101",
		764 =>	x"01010202",
		765 =>	x"02010101",
		766 =>	x"01010101",
		767 =>	x"01010101",
		768 =>	x"01010101", -- IMG_8x8_33_NUM_2
		769 =>	x"01010101",
		770 =>	x"01010102",
		771 =>	x"02010101",
		772 =>	x"01010201",
		773 =>	x"01020101",
		774 =>	x"01010101",
		775 =>	x"01020101",
		776 =>	x"01010102",
		777 =>	x"02010101",
		778 =>	x"01010201",
		779 =>	x"01010101",
		780 =>	x"01010202",
		781 =>	x"02020101",
		782 =>	x"01010101",
		783 =>	x"01010101",
		784 =>	x"01010101", -- IMG_8x8_34_NUM_3
		785 =>	x"01010101",
		786 =>	x"01010202",
		787 =>	x"02010101",
		788 =>	x"01010101",
		789 =>	x"01020101",
		790 =>	x"01010101",
		791 =>	x"02010101",
		792 =>	x"01010101",
		793 =>	x"01020101",
		794 =>	x"01010201",
		795 =>	x"01020101",
		796 =>	x"01010102",
		797 =>	x"02010101",
		798 =>	x"01010101",
		799 =>	x"01010101",
		800 =>	x"01010101", -- IMG_8x8_35_NUM_4
		801 =>	x"01010101",
		802 =>	x"01010201",
		803 =>	x"01010101",
		804 =>	x"01010201",
		805 =>	x"02010101",
		806 =>	x"01010201",
		807 =>	x"02010101",
		808 =>	x"01010202",
		809 =>	x"02020101",
		810 =>	x"01010101",
		811 =>	x"02010101",
		812 =>	x"01010101",
		813 =>	x"02010101",
		814 =>	x"01010101",
		815 =>	x"01010101",
		816 =>	x"01010101", -- IMG_8x8_36_NUM_5
		817 =>	x"01010101",
		818 =>	x"01010202",
		819 =>	x"02020101",
		820 =>	x"01010201",
		821 =>	x"01010101",
		822 =>	x"01010202",
		823 =>	x"02010101",
		824 =>	x"01010101",
		825 =>	x"01020101",
		826 =>	x"01010101",
		827 =>	x"01020101",
		828 =>	x"01010202",
		829 =>	x"02010101",
		830 =>	x"01010101",
		831 =>	x"01010101",
		832 =>	x"01010101", -- IMG_8x8_37_NUM_6
		833 =>	x"01010101",
		834 =>	x"01010102",
		835 =>	x"02020101",
		836 =>	x"01010201",
		837 =>	x"01010101",
		838 =>	x"01010202",
		839 =>	x"02010101",
		840 =>	x"01010201",
		841 =>	x"01020101",
		842 =>	x"01010201",
		843 =>	x"01020101",
		844 =>	x"01010102",
		845 =>	x"02010101",
		846 =>	x"01010101",
		847 =>	x"01010101",
		848 =>	x"01010101", -- IMG_8x8_38_NUM_7
		849 =>	x"01010101",
		850 =>	x"01010202",
		851 =>	x"02020101",
		852 =>	x"01010101",
		853 =>	x"01020101",
		854 =>	x"01010101",
		855 =>	x"02010101",
		856 =>	x"01010102",
		857 =>	x"01010101",
		858 =>	x"01010102",
		859 =>	x"01010101",
		860 =>	x"01010102",
		861 =>	x"01010101",
		862 =>	x"01010101",
		863 =>	x"01010101",
		864 =>	x"01010101", -- IMG_8x8_39_NUM_8
		865 =>	x"01010101",
		866 =>	x"01010102",
		867 =>	x"02010101",
		868 =>	x"01010201",
		869 =>	x"01020101",
		870 =>	x"01010201",
		871 =>	x"01020101",
		872 =>	x"01010102",
		873 =>	x"02010101",
		874 =>	x"01010201",
		875 =>	x"01020101",
		876 =>	x"01010102",
		877 =>	x"02010101",
		878 =>	x"01010101",
		879 =>	x"01010101",
		880 =>	x"01010101", -- IMG_8x8_40_NUM_9
		881 =>	x"01010101",
		882 =>	x"01010102",
		883 =>	x"02010101",
		884 =>	x"01010201",
		885 =>	x"01020101",
		886 =>	x"01010201",
		887 =>	x"01020101",
		888 =>	x"01010102",
		889 =>	x"02020101",
		890 =>	x"01010101",
		891 =>	x"01020101",
		892 =>	x"01010202",
		893 =>	x"02010101",
		894 =>	x"01010101",
		895 =>	x"01010101",
		896 =>	x"01010101", -- IMG_8x8_41_DOTS
		897 =>	x"01010101",
		898 =>	x"01010101",
		899 =>	x"01010101",
		900 =>	x"01010102",
		901 =>	x"01010101",
		902 =>	x"01010101",
		903 =>	x"01010101",
		904 =>	x"01010101",
		905 =>	x"01010101",
		906 =>	x"01010102",
		907 =>	x"01010101",
		908 =>	x"01010101",
		909 =>	x"01010101",
		910 =>	x"01010101",
		911 =>	x"01010101",
		912 =>	x"01010101", -- IMG_8x8_42_FULLSTOP
		913 =>	x"01010101",
		914 =>	x"01010101",
		915 =>	x"01010101",
		916 =>	x"01010101",
		917 =>	x"01010101",
		918 =>	x"01010101",
		919 =>	x"01010101",
		920 =>	x"01010101",
		921 =>	x"01010101",
		922 =>	x"01010102",
		923 =>	x"01010101",
		924 =>	x"01010101",
		925 =>	x"01010101",
		926 =>	x"01010101",
		927 =>	x"01010101",
		928 =>	x"01010101", -- IMG_8x8_BLANK
		929 =>	x"01010101",
		930 =>	x"01010101",
		931 =>	x"01010101",
		932 =>	x"01010101",
		933 =>	x"01010101",
		934 =>	x"01010101",
		935 =>	x"01010101",
		936 =>	x"01010101",
		937 =>	x"01010101",
		938 =>	x"01010101",
		939 =>	x"01010101",
		940 =>	x"01010101",
		941 =>	x"01010101",
		942 =>	x"01010101",
		943 =>	x"01010101",
		944 =>	x"03030303", -- IMG_8x8_BRICK
		945 =>	x"04030303",
		946 =>	x"05050505",
		947 =>	x"04030505",
		948 =>	x"05050505",
		949 =>	x"04030505",
		950 =>	x"04040404",
		951 =>	x"04040404",
		952 =>	x"04030303",
		953 =>	x"03030303",
		954 =>	x"04030505",
		955 =>	x"05050505",
		956 =>	x"04030505",
		957 =>	x"05050505",
		958 =>	x"04040404",
		959 =>	x"04040404",
		960 =>	x"00060606", -- IMG_8x8_GRASS
		961 =>	x"07060800",
		962 =>	x"06060708",
		963 =>	x"06080608",
		964 =>	x"06060606",
		965 =>	x"06080808",
		966 =>	x"07060608",
		967 =>	x"08070608",
		968 =>	x"06060807",
		969 =>	x"08080807",
		970 =>	x"06070608",
		971 =>	x"08080808",
		972 =>	x"08080808",
		973 =>	x"08070808",
		974 =>	x"00080807",
		975 =>	x"08080800",
		976 =>	x"04090902", -- IMG_8x8_ICE
		977 =>	x"04090902",
		978 =>	x"09090909",
		979 =>	x"09090204",
		980 =>	x"09090909",
		981 =>	x"09020409",
		982 =>	x"02090909",
		983 =>	x"02040909",
		984 =>	x"04090902",
		985 =>	x"04090902",
		986 =>	x"09090204",
		987 =>	x"09090204",
		988 =>	x"09020409",
		989 =>	x"09020409",
		990 =>	x"02040909",
		991 =>	x"02040909",
		992 =>	x"09090909", -- IMG_8x8_IRON
		993 =>	x"09090909",
		994 =>	x"09090909",
		995 =>	x"09090904",
		996 =>	x"09090202",
		997 =>	x"02020404",
		998 =>	x"09090202",
		999 =>	x"02020404",
		1000 =>	x"09090202",
		1001 =>	x"02020404",
		1002 =>	x"09090202",
		1003 =>	x"02020404",
		1004 =>	x"09090404",
		1005 =>	x"04040404",
		1006 =>	x"09040404",
		1007 =>	x"04040404",
		1008 =>	x"04040405", -- IMG_8x8_LIVES_REMAINING_ICON
		1009 =>	x"05050404",
		1010 =>	x"04050404",
		1011 =>	x"05040405",
		1012 =>	x"04050405",
		1013 =>	x"05050405",
		1014 =>	x"04050505",
		1015 =>	x"04050505",
		1016 =>	x"04050504",
		1017 =>	x"04040505",
		1018 =>	x"04050505",
		1019 =>	x"04050505",
		1020 =>	x"04050405",
		1021 =>	x"05050405",
		1022 =>	x"04050404",
		1023 =>	x"05040405",
		1024 =>	x"00000000", -- IMG_8x8_NULL
		1025 =>	x"00000000",
		1026 =>	x"00000000",
		1027 =>	x"00000000",
		1028 =>	x"00000000",
		1029 =>	x"00000000",
		1030 =>	x"00000000",
		1031 =>	x"00000000",
		1032 =>	x"00000000",
		1033 =>	x"00000000",
		1034 =>	x"00000000",
		1035 =>	x"00000000",
		1036 =>	x"00000000",
		1037 =>	x"00000000",
		1038 =>	x"00000000",
		1039 =>	x"00000000",
		1040 =>	x"04040404", -- IMG_8x8_TANKS_REMAINING_ICON
		1041 =>	x"04040404",
		1042 =>	x"04000404",
		1043 =>	x"00040400",
		1044 =>	x"04000400",
		1045 =>	x"00000400",
		1046 =>	x"04000000",
		1047 =>	x"03000000",
		1048 =>	x"04000000",
		1049 =>	x"03000000",
		1050 =>	x"04000400",
		1051 =>	x"00000400",
		1052 =>	x"04000404",
		1053 =>	x"00040400",
		1054 =>	x"04040400",
		1055 =>	x"00000404",
		1056 =>	x"0A0A0A0A", -- IMG_8x8_WATER
		1057 =>	x"0A0A0A0B",
		1058 =>	x"0A0B0A0A",
		1059 =>	x"0A0A0A0A",
		1060 =>	x"0A0A0B0A",
		1061 =>	x"0A0A0A0A",
		1062 =>	x"0A0A0A0B",
		1063 =>	x"0A0A0B0A",
		1064 =>	x"0A0A0A0A",
		1065 =>	x"0A0A0A0B",
		1066 =>	x"0A0A0A0B",
		1067 =>	x"0A0A0A0A",
		1068 =>	x"0A0A0B0A",
		1069 =>	x"0B0A0A0A",
		1070 =>	x"0B0A0A0A",
		1071 =>	x"0A0A0A0A",


--			***** 16x16 IMAGES *****


		1072 =>	x"00000000", -- IMG_16x16_BASE_ALIVE
		1073 =>	x"00000000",
		1074 =>	x"00000000",
		1075 =>	x"00000000",
		1076 =>	x"04040000",
		1077 =>	x"00000000",
		1078 =>	x"00000000",
		1079 =>	x"00000404",
		1080 =>	x"00040400",
		1081 =>	x"00000404",
		1082 =>	x"04000000",
		1083 =>	x"00040400",
		1084 =>	x"04040404",
		1085 =>	x"00000004",
		1086 =>	x"03040000",
		1087 =>	x"04040404",
		1088 =>	x"00040404",
		1089 =>	x"00000004",
		1090 =>	x"04000000",
		1091 =>	x"04040400",
		1092 =>	x"04040404",
		1093 =>	x"04040004",
		1094 =>	x"04000404",
		1095 =>	x"04040404",
		1096 =>	x"00000403",
		1097 =>	x"04040404",
		1098 =>	x"04040404",
		1099 =>	x"03040000",
		1100 =>	x"00040404",
		1101 =>	x"03040404",
		1102 =>	x"04040403",
		1103 =>	x"04040400",
		1104 =>	x"00000404",
		1105 =>	x"04040304",
		1106 =>	x"04030404",
		1107 =>	x"04040000",
		1108 =>	x"00000404",
		1109 =>	x"04040404",
		1110 =>	x"04040404",
		1111 =>	x"04040000",
		1112 =>	x"00000004",
		1113 =>	x"04040004",
		1114 =>	x"04000404",
		1115 =>	x"04000000",
		1116 =>	x"00000000",
		1117 =>	x"00000004",
		1118 =>	x"04000000",
		1119 =>	x"00000000",
		1120 =>	x"00000000",
		1121 =>	x"00000404",
		1122 =>	x"04040000",
		1123 =>	x"00000000",
		1124 =>	x"00000000",
		1125 =>	x"04040404",
		1126 =>	x"04040404",
		1127 =>	x"00000000",
		1128 =>	x"00000000",
		1129 =>	x"04040004",
		1130 =>	x"04000404",
		1131 =>	x"00000000",
		1132 =>	x"00000000",
		1133 =>	x"00000000",
		1134 =>	x"00000000",
		1135 =>	x"00000000",
		1136 =>	x"00000000", -- IMG_16x16_BASE_DEAD
		1137 =>	x"00000000",
		1138 =>	x"00000000",
		1139 =>	x"00000000",
		1140 =>	x"00000000",
		1141 =>	x"00050000",
		1142 =>	x"00000000",
		1143 =>	x"00000000",
		1144 =>	x"00000000",
		1145 =>	x"05050004",
		1146 =>	x"00000000",
		1147 =>	x"00000000",
		1148 =>	x"00000000",
		1149 =>	x"05000404",
		1150 =>	x"04000000",
		1151 =>	x"00000000",
		1152 =>	x"00000005",
		1153 =>	x"00040404",
		1154 =>	x"04040000",
		1155 =>	x"00000000",
		1156 =>	x"00000505",
		1157 =>	x"00040404",
		1158 =>	x"04040404",
		1159 =>	x"04000000",
		1160 =>	x"00000500",
		1161 =>	x"04040404",
		1162 =>	x"04040404",
		1163 =>	x"04040000",
		1164 =>	x"00050500",
		1165 =>	x"04040404",
		1166 =>	x"04040404",
		1167 =>	x"04040000",
		1168 =>	x"00050000",
		1169 =>	x"04040404",
		1170 =>	x"04040404",
		1171 =>	x"00040400",
		1172 =>	x"00050004",
		1173 =>	x"04040404",
		1174 =>	x"04000004",
		1175 =>	x"00040400",
		1176 =>	x"00050000",
		1177 =>	x"00040404",
		1178 =>	x"00000000",
		1179 =>	x"00040000",
		1180 =>	x"00050000",
		1181 =>	x"00000004",
		1182 =>	x"00000000",
		1183 =>	x"00040000",
		1184 =>	x"00050000",
		1185 =>	x"00000000",
		1186 =>	x"00000000",
		1187 =>	x"00000000",
		1188 =>	x"00050000",
		1189 =>	x"00000000",
		1190 =>	x"00000000",
		1191 =>	x"00000000",
		1192 =>	x"00050000",
		1193 =>	x"00000000",
		1194 =>	x"00000000",
		1195 =>	x"00000000",
		1196 =>	x"00000000",
		1197 =>	x"00000000",
		1198 =>	x"00000000",
		1199 =>	x"00000000",
		1200 =>	x"00000000", -- IMG_16x16_BONUS_BOMB
		1201 =>	x"00000000",
		1202 =>	x"00000000",
		1203 =>	x"00000000",
		1204 =>	x"00020202",
		1205 =>	x"02020202",
		1206 =>	x"02020202",
		1207 =>	x"02020900",
		1208 =>	x"02000000",
		1209 =>	x"00000000",
		1210 =>	x"00000000",
		1211 =>	x"0000020C",
		1212 =>	x"02000C0C",
		1213 =>	x"0C020202",
		1214 =>	x"0909000C",
		1215 =>	x"0C0C020C",
		1216 =>	x"02000C0C",
		1217 =>	x"0C02090C",
		1218 =>	x"00000900",
		1219 =>	x"0C0C020C",
		1220 =>	x"02000C0C",
		1221 =>	x"02090909",
		1222 =>	x"0C000009",
		1223 =>	x"000C020C",
		1224 =>	x"02000C02",
		1225 =>	x"090C0209",
		1226 =>	x"0C090009",
		1227 =>	x"000C020C",
		1228 =>	x"02000C09",
		1229 =>	x"00090000",
		1230 =>	x"09000009",
		1231 =>	x"000C020C",
		1232 =>	x"02000C02",
		1233 =>	x"090C0209",
		1234 =>	x"0C090009",
		1235 =>	x"000C020C",
		1236 =>	x"02000C09",
		1237 =>	x"00090000",
		1238 =>	x"09000009",
		1239 =>	x"000C020C",
		1240 =>	x"02000C02",
		1241 =>	x"090C0209",
		1242 =>	x"0C090000",
		1243 =>	x"0C0C020C",
		1244 =>	x"02000C0C",
		1245 =>	x"090C0000",
		1246 =>	x"09000C0C",
		1247 =>	x"0C0C020C",
		1248 =>	x"02000C0C",
		1249 =>	x"0C020909",
		1250 =>	x"000C0C0C",
		1251 =>	x"0C0C020C",
		1252 =>	x"02000C0C",
		1253 =>	x"0C000000",
		1254 =>	x"0C0C0C0C",
		1255 =>	x"0C0C020C",
		1256 =>	x"09020202",
		1257 =>	x"02020202",
		1258 =>	x"02020202",
		1259 =>	x"0202090C",
		1260 =>	x"000C0C0C",
		1261 =>	x"0C0C0C0C",
		1262 =>	x"0C0C0C0C",
		1263 =>	x"0C0C0C00",
		1264 => x"02020202", -- IMG_16x16_MAIN_TANK_B
		1265 => x"02020202",
		1266 => x"1F1F1F1F",
		1267 => x"1F1F1F1F",
		1268 => x"1F1F1F1F",
		1269 => x"1F1F1F1F",
		1270 => x"1F1F1F1F",
		1271 => x"1F1F1F1F",
		1272 => x"1F1F1F1F",
		1273 => x"1F1F1F0F",
		1274 => x"1F1F1F1F",
		1275 => x"1F1F1F1F",
		1276 => x"1F1F1F1F",
		1277 => x"1F1F1F0F",
		1278 => x"1F1F1F1F",
		1279 => x"1F1F1F1F",
		1280 => x"1F111110",
		1281 => x"1F1F1F0F",
		1282 => x"1F1F1F0F",
		1283 => x"11111F1F",
		1284 => x"1F0F100F",
		1285 => x"1F1F1F0F",
		1286 => x"1F1F1F11",
		1287 => x"10101F1F",
		1288 => x"1F11110F",
		1289 => x"1F0F100F",
		1290 => x"11111F11",
		1291 => x"11111F1F",
		1292 => x"1F0F100F",
		1293 => x"0F0F1010",
		1294 => x"10101111",
		1295 => x"10101F1F",
		1296 => x"1F11110F",
		1297 => x"0F100F0F",
		1298 => x"10101011",
		1299 => x"11111F1F",
		1300 => x"1F0F100F",
		1301 => x"0F100F10",
		1302 => x"11101011",
		1303 => x"10101F1F",
		1304 => x"1F11110F",
		1305 => x"0F100F10",
		1306 => x"11101011",
		1307 => x"11111F1F",
		1308 => x"1F0F100F",
		1309 => x"0F0F1011",
		1310 => x"11101011",
		1311 => x"10101F1F",
		1312 => x"1F11110F",
		1313 => x"110F0F10",
		1314 => x"10101111",
		1315 => x"11111F1F",
		1316 => x"1F0F100F",
		1317 => x"1F111111",
		1318 => x"11111F11",
		1319 => x"10101F1F",
		1320 => x"1F111110",
		1321 => x"1F1F1F1F",
		1322 => x"1F1F1F11",
		1323 => x"11111F1F",
		1324 => x"1F1F1F1F",
		1325 => x"1F1F1F1F",
		1326 => x"1F1F1F1F",
		1327 => x"1F1F1F1F",
		1328 => x"1F1F1F1F", -- IMG_16x16_ENEMY_TANK1_B
		1329 => x"1F1F1F1F",
		1330 => x"1F1F1F1F",
		1331 => x"1F1F1F1F",
		1332 => x"1F1F1F1F",
		1333 => x"1F1F1F02",
		1334 => x"1F1F1F1F",
		1335 => x"1F1F1F1F",
		1336 => x"1F1F1F1F",
		1337 => x"1F1F1F02",
		1338 => x"1F1F1F1F",
		1339 => x"1F1F1F1F",
		1340 => x"1F1F1F1F",
		1341 => x"1F1F1F02",
		1342 => x"1F1F1F1F",
		1343 => x"1F1F1F1F",
		1344 => x"1F0C0C09",
		1345 => x"1F1F0902",
		1346 => x"0C1F1F02",
		1347 => x"0C0C1F1F",
		1348 => x"1F020909",
		1349 => x"1F020902",
		1350 => x"0C0C1F09",
		1351 => x"09091F1F",
		1352 => x"1F0C0C09",
		1353 => x"02020902",
		1354 => x"0C0C0C09",
		1355 => x"0C0C1F1F",
		1356 => x"1F020909",
		1357 => x"02020909",
		1358 => x"090C0C09",
		1359 => x"09091F1F",
		1360 => x"1F0C0C09",
		1361 => x"0209090C",
		1362 => x"09090C09",
		1363 => x"0C0C1F1F",
		1364 => x"1F020909",
		1365 => x"02090C0C",
		1366 => x"02090C09",
		1367 => x"09091F1F",
		1368 => x"1F0C0C09",
		1369 => x"02090C02",
		1370 => x"02090C09",
		1371 => x"0C0C1F1F",
		1372 => x"1F020909",
		1373 => x"02090909",
		1374 => x"09090C09",
		1375 => x"09091F1F",
		1376 => x"1F0C0C09",
		1377 => x"02020909",
		1378 => x"090C0C09",
		1379 => x"0C0C1F1F",
		1380 => x"1F020909",
		1381 => x"1F020909",
		1382 => x"0C0C1F09",
		1383 => x"09091F1F",
		1384 => x"1F0C0C09",
		1385 => x"1F1F0C0C",
		1386 => x"0C1F1F09",
		1387 => x"0C0C1F1F",
		1388 => x"1F1F1F1F",
		1389 => x"1F1F1F09",
		1390 => x"1F1F1F1F",
		1391 => x"1F1F1F1F",
		1392 =>	x"00000000", -- IMG_16x16_BONUS_SHOVEL
		1393 =>	x"00000000",
		1394 =>	x"00000000",
		1395 =>	x"00000000",
		1396 =>	x"00020202",
		1397 =>	x"02020202",
		1398 =>	x"02020202",
		1399 =>	x"02020900",
		1400 =>	x"02000000",
		1401 =>	x"00000000",
		1402 =>	x"00000000",
		1403 =>	x"0000020C",
		1404 =>	x"02000C0C",
		1405 =>	x"0C0C0C0C",
		1406 =>	x"0C0C020C",
		1407 =>	x"0C0C020C",
		1408 =>	x"02000C0C",
		1409 =>	x"0C0C0C0C",
		1410 =>	x"0C0C0209",
		1411 =>	x"0C0C020C",
		1412 =>	x"02000C0C",
		1413 =>	x"0C0C0C0C",
		1414 =>	x"0C0C0909",
		1415 =>	x"090C020C",
		1416 =>	x"02000C0C",
		1417 =>	x"0C0C0C0C",
		1418 =>	x"0C020000",
		1419 =>	x"000C020C",
		1420 =>	x"02000C0C",
		1421 =>	x"0C020C0C",
		1422 =>	x"02000C0C",
		1423 =>	x"0C0C020C",
		1424 =>	x"02000C0C",
		1425 =>	x"02020902",
		1426 =>	x"000C0C0C",
		1427 =>	x"0C0C020C",
		1428 =>	x"02000C02",
		1429 =>	x"02090C09",
		1430 =>	x"000C0C0C",
		1431 =>	x"0C0C020C",
		1432 =>	x"02000C02",
		1433 =>	x"090C0909",
		1434 =>	x"09000C0C",
		1435 =>	x"0C0C020C",
		1436 =>	x"02000C09",
		1437 =>	x"09090909",
		1438 =>	x"000C0C0C",
		1439 =>	x"0C0C020C",
		1440 =>	x"02000C09",
		1441 =>	x"09090900",
		1442 =>	x"0C0C0C0C",
		1443 =>	x"0C0C020C",
		1444 =>	x"02000C00",
		1445 =>	x"0000000C",
		1446 =>	x"0C0C0C0C",
		1447 =>	x"0C0C020C",
		1448 =>	x"09020202",
		1449 =>	x"02020202",
		1450 =>	x"02020202",
		1451 =>	x"0202090C",
		1452 =>	x"000C0C0C",
		1453 =>	x"0C0C0C0C",
		1454 =>	x"0C0C0C0C",
		1455 =>	x"0C0C0C00",
		1456 =>	x"00000000", -- IMG_16x16_BONUS_STAR
		1457 =>	x"00000000",
		1458 =>	x"00000000",
		1459 =>	x"00000000",
		1460 =>	x"00020202",
		1461 =>	x"02020202",
		1462 =>	x"02020202",
		1463 =>	x"02020900",
		1464 =>	x"02000000",
		1465 =>	x"00000000",
		1466 =>	x"00000000",
		1467 =>	x"0000020C",
		1468 =>	x"02000C0C",
		1469 =>	x"0C0C0C02",
		1470 =>	x"000C0C0C",
		1471 =>	x"0C0C020C",
		1472 =>	x"02000C0C",
		1473 =>	x"0C0C0202",
		1474 =>	x"09000C0C",
		1475 =>	x"0C0C020C",
		1476 =>	x"02000C0C",
		1477 =>	x"0C0C0202",
		1478 =>	x"09000C0C",
		1479 =>	x"0C0C020C",
		1480 =>	x"02000202",
		1481 =>	x"02020209",
		1482 =>	x"09020202",
		1483 =>	x"0200020C",
		1484 =>	x"02000C09",
		1485 =>	x"09090209",
		1486 =>	x"02090909",
		1487 =>	x"0000020C",
		1488 =>	x"02000C0C",
		1489 =>	x"09020202",
		1490 =>	x"02090900",
		1491 =>	x"000C020C",
		1492 =>	x"02000C0C",
		1493 =>	x"02020909",
		1494 =>	x"02020900",
		1495 =>	x"0C0C020C",
		1496 =>	x"02000C09",
		1497 =>	x"02090900",
		1498 =>	x"09090209",
		1499 =>	x"000C020C",
		1500 =>	x"02000C02",
		1501 =>	x"09090000",
		1502 =>	x"00090902",
		1503 =>	x"000C020C",
		1504 =>	x"02000C09",
		1505 =>	x"0000000C",
		1506 =>	x"0C000009",
		1507 =>	x"000C020C",
		1508 =>	x"02000C00",
		1509 =>	x"000C0C0C",
		1510 =>	x"0C0C0C00",
		1511 =>	x"000C020C",
		1512 =>	x"09020202",
		1513 =>	x"02020202",
		1514 =>	x"02020202",
		1515 =>	x"0202090C",
		1516 =>	x"000C0C0C",
		1517 =>	x"0C0C0C0C",
		1518 =>	x"0C0C0C0C",
		1519 =>	x"0C0C0C00",
		1520 =>	x"00000000", -- IMG_16x16_BONUS_TANK
		1521 =>	x"00000000",
		1522 =>	x"00000000",
		1523 =>	x"00000000",
		1524 =>	x"00020202",
		1525 =>	x"02020202",
		1526 =>	x"02020202",
		1527 =>	x"02020900",
		1528 =>	x"02000000",
		1529 =>	x"00000000",
		1530 =>	x"00000000",
		1531 =>	x"0000020C",
		1532 =>	x"02000C0C",
		1533 =>	x"0C0C0C0C",
		1534 =>	x"0C0C0C0C",
		1535 =>	x"0C0C020C",
		1536 =>	x"02000C02",
		1537 =>	x"0C0C0C0C",
		1538 =>	x"0C0C0C0C",
		1539 =>	x"0C0C020C",
		1540 =>	x"02000902",
		1541 =>	x"02020202",
		1542 =>	x"02020900",
		1543 =>	x"0C0C020C",
		1544 =>	x"02000209",
		1545 =>	x"09090909",
		1546 =>	x"09090909",
		1547 =>	x"000C020C",
		1548 =>	x"02000009",
		1549 =>	x"090C0C0C",
		1550 =>	x"0C0C0C09",
		1551 =>	x"000C020C",
		1552 =>	x"02000C00",
		1553 =>	x"0009090C",
		1554 =>	x"09090909",
		1555 =>	x"0900020C",
		1556 =>	x"02000C0C",
		1557 =>	x"0C000900",
		1558 =>	x"0009020C",
		1559 =>	x"0900020C",
		1560 =>	x"02000C0C",
		1561 =>	x"0C0C0009",
		1562 =>	x"0909020C",
		1563 =>	x"0900020C",
		1564 =>	x"02000C0C",
		1565 =>	x"0C0C0C00",
		1566 =>	x"00090C0C",
		1567 =>	x"0900020C",
		1568 =>	x"02000C0C",
		1569 =>	x"0C0C0C0C",
		1570 =>	x"0C090909",
		1571 =>	x"0900020C",
		1572 =>	x"02000C0C",
		1573 =>	x"0C0C0C0C",
		1574 =>	x"0C000000",
		1575 =>	x"000C020C",
		1576 =>	x"09020202",
		1577 =>	x"02020202",
		1578 =>	x"02020202",
		1579 =>	x"0202090C",
		1580 =>	x"000C0C0C",
		1581 =>	x"0C0C0C0C",
		1582 =>	x"0C0C0C0C",
		1583 =>	x"0C0C0C00",
		1584 =>	x"00000000", -- IMG_16x16_BONUS_TIME
		1585 =>	x"00000000",
		1586 =>	x"00000000",
		1587 =>	x"00000000",
		1588 =>	x"00000202",
		1589 =>	x"02020202",
		1590 =>	x"02020202",
		1591 =>	x"02020209",
		1592 =>	x"0C020000",
		1593 =>	x"00000000",
		1594 =>	x"00000000",
		1595 =>	x"00000002",
		1596 =>	x"0C02000C",
		1597 =>	x"0C0C0C02",
		1598 =>	x"09020900",
		1599 =>	x"0C0C0C02",
		1600 =>	x"0C02000C",
		1601 =>	x"0C0C0C09",
		1602 =>	x"00000002",
		1603 =>	x"09000C02",
		1604 =>	x"0C02000C",
		1605 =>	x"0C0C0909",
		1606 =>	x"09090000",
		1607 =>	x"00000C02",
		1608 =>	x"0C02000C",
		1609 =>	x"0C090202",
		1610 =>	x"02020900",
		1611 =>	x"0C0C0C02",
		1612 =>	x"0C02000C",
		1613 =>	x"0902020C",
		1614 =>	x"02020209",
		1615 =>	x"000C0C02",
		1616 =>	x"0C02000C",
		1617 =>	x"0902020C",
		1618 =>	x"02020209",
		1619 =>	x"000C0C02",
		1620 =>	x"0C02000C",
		1621 =>	x"09020202",
		1622 =>	x"0C020209",
		1623 =>	x"000C0C02",
		1624 =>	x"0C02000C",
		1625 =>	x"00090202",
		1626 =>	x"02020900",
		1627 =>	x"0C0C0C02",
		1628 =>	x"0C02000C",
		1629 =>	x"0C000909",
		1630 =>	x"0909000C",
		1631 =>	x"0C0C0C02",
		1632 =>	x"0C02000C",
		1633 =>	x"0C0C0000",
		1634 =>	x"00000C0C",
		1635 =>	x"0C0C0C02",
		1636 =>	x"0C02000C",
		1637 =>	x"0C0C0C0C",
		1638 =>	x"0C0C0C0C",
		1639 =>	x"0C0C0C02",
		1640 =>	x"0C090202",
		1641 =>	x"02020202",
		1642 =>	x"02020202",
		1643 =>	x"02020209",
		1644 =>	x"00000C0C",
		1645 =>	x"0C0C0C0C",
		1646 =>	x"0C0C0C0C",
		1647 =>	x"0C0C0C0C",
		1648 =>	x"00000000", -- IMG_16x16_BULLET
		1649 =>	x"00000000",
		1650 =>	x"00000000",
		1651 =>	x"00000000",
		1652 =>	x"00000000",
		1653 =>	x"00000000",
		1654 =>	x"00000000",
		1655 =>	x"00000000",
		1656 =>	x"00000000",
		1657 =>	x"00000000",
		1658 =>	x"00000000",
		1659 =>	x"00000000",
		1660 =>	x"00000000",
		1661 =>	x"00000000",
		1662 =>	x"00000000",
		1663 =>	x"00000000",
		1664 =>	x"00000000",
		1665 =>	x"00000000",
		1666 =>	x"00000000",
		1667 =>	x"00000000",
		1668 =>	x"00000000",
		1669 =>	x"00000009",
		1670 =>	x"00000000",
		1671 =>	x"00000000",
		1672 =>	x"00000000",
		1673 =>	x"00000909",
		1674 =>	x"09000000",
		1675 =>	x"00000000",
		1676 =>	x"00000000",
		1677 =>	x"00000909",
		1678 =>	x"09000000",
		1679 =>	x"00000000",
		1680 =>	x"00000000",
		1681 =>	x"00000909",
		1682 =>	x"09000000",
		1683 =>	x"00000000",
		1684 =>	x"00000000",
		1685 =>	x"00000000",
		1686 =>	x"00000000",
		1687 =>	x"00000000",
		1688 =>	x"00000000",
		1689 =>	x"00000000",
		1690 =>	x"00000000",
		1691 =>	x"00000000",
		1692 =>	x"00000000",
		1693 =>	x"00000000",
		1694 =>	x"00000000",
		1695 =>	x"00000000",
		1696 =>	x"00000000",
		1697 =>	x"00000000",
		1698 =>	x"00000000",
		1699 =>	x"00000000",
		1700 =>	x"00000000",
		1701 =>	x"00000000",
		1702 =>	x"00000000",
		1703 =>	x"00000000",
		1704 =>	x"00000000",
		1705 =>	x"00000000",
		1706 =>	x"00000000",
		1707 =>	x"00000000",
		1708 =>	x"00000000",
		1709 =>	x"00000000",
		1710 =>	x"00000000",
		1711 =>	x"00000000",
		1712 =>	x"00000000", -- IMG_16x16_ENEMY_TANK1
		1713 =>	x"00000000",
		1714 =>	x"00000000",
		1715 =>	x"00000000",
		1716 =>	x"00000000",
		1717 =>	x"00000002",
		1718 =>	x"00000000",
		1719 =>	x"00000000",
		1720 =>	x"00000000",
		1721 =>	x"00000002",
		1722 =>	x"00000000",
		1723 =>	x"00000000",
		1724 =>	x"00000000",
		1725 =>	x"00000002",
		1726 =>	x"00000000",
		1727 =>	x"00000000",
		1728 =>	x"00020909",
		1729 =>	x"00000902",
		1730 =>	x"0C000002",
		1731 =>	x"09090000",
		1732 =>	x"000C0C09",
		1733 =>	x"00020902",
		1734 =>	x"0C0C0009",
		1735 =>	x"0C0C0000",
		1736 =>	x"00020909",
		1737 =>	x"02020902",
		1738 =>	x"0C0C0C09",
		1739 =>	x"09090000",
		1740 =>	x"000C0C09",
		1741 =>	x"02020909",
		1742 =>	x"090C0C09",
		1743 =>	x"0C0C0000",
		1744 =>	x"00020909",
		1745 =>	x"0209090C",
		1746 =>	x"09090C09",
		1747 =>	x"09090000",
		1748 =>	x"000C0C09",
		1749 =>	x"02090C0C",
		1750 =>	x"02090C09",
		1751 =>	x"0C0C0000",
		1752 =>	x"00020909",
		1753 =>	x"02090C02",
		1754 =>	x"02090C09",
		1755 =>	x"09090000",
		1756 =>	x"000C0C09",
		1757 =>	x"02090909",
		1758 =>	x"09090C09",
		1759 =>	x"0C0C0000",
		1760 =>	x"00020909",
		1761 =>	x"02020909",
		1762 =>	x"090C0C09",
		1763 =>	x"09090000",
		1764 =>	x"000C0C09",
		1765 =>	x"00020909",
		1766 =>	x"0C0C0009",
		1767 =>	x"0C0C0000",
		1768 =>	x"00020909",
		1769 =>	x"00000C0C",
		1770 =>	x"0C000009",
		1771 =>	x"09090000",
		1772 =>	x"00000000",
		1773 =>	x"00000009",
		1774 =>	x"00000000",
		1775 =>	x"00000000",
		1776 =>	x"00000000", -- IMG_16x16_ENEMY_TANK2
		1777 =>	x"00000000",
		1778 =>	x"00000000",
		1779 =>	x"00000000",
		1780 =>	x"00000000",
		1781 =>	x"00000002",
		1782 =>	x"00000000",
		1783 =>	x"00000000",
		1784 =>	x"00000000",
		1785 =>	x"00000002",
		1786 =>	x"00000000",
		1787 =>	x"00000000",
		1788 =>	x"00090C00",
		1789 =>	x"02020C02",
		1790 =>	x"0C090900",
		1791 =>	x"090C0000",
		1792 =>	x"000C0C02",
		1793 =>	x"02020C02",
		1794 =>	x"0C090909",
		1795 =>	x"0C0C0000",
		1796 =>	x"000C0C09",
		1797 =>	x"02020C02",
		1798 =>	x"0C0C0C09",
		1799 =>	x"0C0C0000",
		1800 =>	x"00000009",
		1801 =>	x"09020902",
		1802 =>	x"090C0C09",
		1803 =>	x"00000000",
		1804 =>	x"00000009",
		1805 =>	x"02090909",
		1806 =>	x"09090C09",
		1807 =>	x"00000000",
		1808 =>	x"00090C09",
		1809 =>	x"0209090C",
		1810 =>	x"09090C09",
		1811 =>	x"090C0000",
		1812 =>	x"000C0C09",
		1813 =>	x"02090C0C",
		1814 =>	x"02090C09",
		1815 =>	x"0C0C0000",
		1816 =>	x"000C0C09",
		1817 =>	x"02090C02",
		1818 =>	x"02090C09",
		1819 =>	x"0C0C0000",
		1820 =>	x"00000009",
		1821 =>	x"02090909",
		1822 =>	x"09090C09",
		1823 =>	x"00000000",
		1824 =>	x"00000009",
		1825 =>	x"02020909",
		1826 =>	x"09020C09",
		1827 =>	x"00000000",
		1828 =>	x"00090C09",
		1829 =>	x"09090202",
		1830 =>	x"020C0C09",
		1831 =>	x"090C0000",
		1832 =>	x"000C0C09",
		1833 =>	x"0C0C0C0C",
		1834 =>	x"0C0C0C09",
		1835 =>	x"0C0C0000",
		1836 =>	x"000C0C00",
		1837 =>	x"0C0C0C02",
		1838 =>	x"0C0C0C00",
		1839 =>	x"0C0C0000",
		1840 =>	x"00000000", -- IMG_16x16_ENEMY_TANK3
		1841 =>	x"00000000",
		1842 =>	x"00000000",
		1843 =>	x"00000000",
		1844 =>	x"00000000",
		1845 =>	x"00000202",
		1846 =>	x"09000000",
		1847 =>	x"00000000",
		1848 =>	x"00000000",
		1849 =>	x"00000002",
		1850 =>	x"00000000",
		1851 =>	x"00000000",
		1852 =>	x"00000000",
		1853 =>	x"00000002",
		1854 =>	x"00000000",
		1855 =>	x"00000000",
		1856 =>	x"00020909",
		1857 =>	x"00000902",
		1858 =>	x"0C000002",
		1859 =>	x"09090000",
		1860 =>	x"000C0C09",
		1861 =>	x"00020902",
		1862 =>	x"0C0C0009",
		1863 =>	x"0C0C0000",
		1864 =>	x"00020909",
		1865 =>	x"02020902",
		1866 =>	x"0C0C0C09",
		1867 =>	x"09090000",
		1868 =>	x"000C0C09",
		1869 =>	x"02020909",
		1870 =>	x"090C0C09",
		1871 =>	x"0C0C0000",
		1872 =>	x"00020909",
		1873 =>	x"0209090C",
		1874 =>	x"09090C09",
		1875 =>	x"09090000",
		1876 =>	x"000C0C09",
		1877 =>	x"02090C0C",
		1878 =>	x"02090C09",
		1879 =>	x"0C0C0000",
		1880 =>	x"00020909",
		1881 =>	x"02090C02",
		1882 =>	x"02090C09",
		1883 =>	x"09090000",
		1884 =>	x"000C0C09",
		1885 =>	x"02090909",
		1886 =>	x"09090C09",
		1887 =>	x"0C0C0000",
		1888 =>	x"00020909",
		1889 =>	x"02020909",
		1890 =>	x"090C0C09",
		1891 =>	x"09090000",
		1892 =>	x"000C0C09",
		1893 =>	x"00020209",
		1894 =>	x"0C0C0009",
		1895 =>	x"0C0C0000",
		1896 =>	x"00020909",
		1897 =>	x"0002020C",
		1898 =>	x"0C0C0009",
		1899 =>	x"09090000",
		1900 =>	x"000C0C09",
		1901 =>	x"00000902",
		1902 =>	x"0C000009",
		1903 =>	x"0C0C0000",
		1904 =>	x"00000000", -- IMG_16x16_ENEMY_TANK4
		1905 =>	x"00000000",
		1906 =>	x"00000000",
		1907 =>	x"00000000",
		1908 =>	x"00020909",
		1909 =>	x"00000202",
		1910 =>	x"09000002",
		1911 =>	x"09090000",
		1912 =>	x"000C0C09",
		1913 =>	x"090C0202",
		1914 =>	x"090C0909",
		1915 =>	x"0C0C0000",
		1916 =>	x"00020909",
		1917 =>	x"09090902",
		1918 =>	x"0C090909",
		1919 =>	x"09090000",
		1920 =>	x"000C0C09",
		1921 =>	x"02090902",
		1922 =>	x"0C09090C",
		1923 =>	x"0C0C0000",
		1924 =>	x"00020909",
		1925 =>	x"02090902",
		1926 =>	x"0C02090C",
		1927 =>	x"09090000",
		1928 =>	x"000C0C09",
		1929 =>	x"02020902",
		1930 =>	x"0C020C0C",
		1931 =>	x"0C0C0000",
		1932 =>	x"00020909",
		1933 =>	x"02020202",
		1934 =>	x"02020C0C",
		1935 =>	x"09090000",
		1936 =>	x"000C0C09",
		1937 =>	x"0209090C",
		1938 =>	x"09090C0C",
		1939 =>	x"0C0C0000",
		1940 =>	x"00020909",
		1941 =>	x"02090C0C",
		1942 =>	x"02090C0C",
		1943 =>	x"09090000",
		1944 =>	x"000C0C09",
		1945 =>	x"02090C02",
		1946 =>	x"02090C0C",
		1947 =>	x"0C0C0000",
		1948 =>	x"00020909",
		1949 =>	x"02090909",
		1950 =>	x"09090C0C",
		1951 =>	x"09090000",
		1952 =>	x"000C0C09",
		1953 =>	x"02090909",
		1954 =>	x"09090C0C",
		1955 =>	x"0C0C0000",
		1956 =>	x"00020909",
		1957 =>	x"090C0C0C",
		1958 =>	x"0C0C090C",
		1959 =>	x"09090000",
		1960 =>	x"000C0C09",
		1961 =>	x"0C0C0C0C",
		1962 =>	x"0C0C0C09",
		1963 =>	x"0C0C0000",
		1964 =>	x"00020909",
		1965 =>	x"00000009",
		1966 =>	x"0000000C",
		1967 =>	x"09090000",
		1968 =>	x"00000000", -- IMG_16x16_EXPLOSION
		1969 =>	x"0D000D00",
		1970 =>	x"0000000D",
		1971 =>	x"00000D00",
		1972 =>	x"00020000",
		1973 =>	x"00020000",
		1974 =>	x"02000D00",
		1975 =>	x"00020D00",
		1976 =>	x"000D0D02",
		1977 =>	x"02000002",
		1978 =>	x"02000000",
		1979 =>	x"020D0000",
		1980 =>	x"00000D0D",
		1981 =>	x"020D0D02",
		1982 =>	x"0D0D0002",
		1983 =>	x"020D0000",
		1984 =>	x"0000000D",
		1985 =>	x"0E020202",
		1986 =>	x"020D0202",
		1987 =>	x"0D0D000D",
		1988 =>	x"0002000D",
		1989 =>	x"02020E02",
		1990 =>	x"0002020E",
		1991 =>	x"0D000000",
		1992 =>	x"00000D02",
		1993 =>	x"020E0D0E",
		1994 =>	x"0E000E0D",
		1995 =>	x"020D0000",
		1996 =>	x"02020202",
		1997 =>	x"00020E00",
		1998 =>	x"000E0202",
		1999 =>	x"02020202",
		2000 =>	x"000D0D0D",
		2001 =>	x"02020D0E",
		2002 =>	x"000E020D",
		2003 =>	x"0D0D0000",
		2004 =>	x"0000000D",
		2005 =>	x"0D0D0002",
		2006 =>	x"0E000D0D",
		2007 =>	x"02020000",
		2008 =>	x"00020D0D",
		2009 =>	x"02020D02",
		2010 =>	x"00020E02",
		2011 =>	x"0D0D0200",
		2012 =>	x"00000202",
		2013 =>	x"020E020D",
		2014 =>	x"020D0202",
		2015 =>	x"00000000",
		2016 =>	x"000D020D",
		2017 =>	x"0D020D02",
		2018 =>	x"020D0D02",
		2019 =>	x"02000D00",
		2020 =>	x"00020D00",
		2021 =>	x"000D000D",
		2022 =>	x"020D000D",
		2023 =>	x"0D020000",
		2024 =>	x"020D0000",
		2025 =>	x"0D000000",
		2026 =>	x"02000000",
		2027 =>	x"000D0200",
		2028 =>	x"00000000",
		2029 =>	x"00000000",
		2030 =>	x"02000D00",
		2031 =>	x"00000D00",
		2032 =>	x"00000404", -- IMG_16x16_FLAG
		2033 =>	x"04040404",
		2034 =>	x"04040404",
		2035 =>	x"04040404",
		2036 =>	x"00000505",
		2037 =>	x"04040404",
		2038 =>	x"04040404",
		2039 =>	x"04040404",
		2040 =>	x"00000505",
		2041 =>	x"05050404",
		2042 =>	x"04040404",
		2043 =>	x"04040404",
		2044 =>	x"00000505",
		2045 =>	x"05050505",
		2046 =>	x"04040404",
		2047 =>	x"04040404",
		2048 =>	x"00000505",
		2049 =>	x"05050505",
		2050 =>	x"05050404",
		2051 =>	x"04040404",
		2052 =>	x"00000505",
		2053 =>	x"05050505",
		2054 =>	x"05050505",
		2055 =>	x"04040404",
		2056 =>	x"00000505",
		2057 =>	x"05050505",
		2058 =>	x"05050505",
		2059 =>	x"05050404",
		2060 =>	x"00000505",
		2061 =>	x"05050505",
		2062 =>	x"05050505",
		2063 =>	x"05050505",
		2064 =>	x"00000505",
		2065 =>	x"05050505",
		2066 =>	x"05050505",
		2067 =>	x"05050505",
		2068 =>	x"00000404",
		2069 =>	x"04040404",
		2070 =>	x"04040404",
		2071 =>	x"04040404",
		2072 =>	x"00000404",
		2073 =>	x"04040404",
		2074 =>	x"04040404",
		2075 =>	x"04040404",
		2076 =>	x"00000404",
		2077 =>	x"04040404",
		2078 =>	x"04040404",
		2079 =>	x"04040404",
		2080 =>	x"00000404",
		2081 =>	x"04040404",
		2082 =>	x"04040404",
		2083 =>	x"04040404",
		2084 =>	x"00000404",
		2085 =>	x"04040404",
		2086 =>	x"04040404",
		2087 =>	x"04040404",
		2088 =>	x"00000404",
		2089 =>	x"04040404",
		2090 =>	x"04040404",
		2091 =>	x"04040404",
		2092 =>	x"04040404",
		2093 =>	x"04040404",
		2094 =>	x"04040404",
		2095 =>	x"04040404",
		2096 =>	x"00000000", -- IMG_16x16_MAIN_TANK
		2097 =>	x"00000000",
		2098 =>	x"00000000",
		2099 =>	x"00000000",
		2100 =>	x"00000000",
		2101 =>	x"00000000",
		2102 =>	x"00000000",
		2103 =>	x"00000000",
		2104 =>	x"00000000",
		2105 =>	x"0000000F",
		2106 =>	x"00000000",
		2107 =>	x"00000000",
		2108 =>	x"00000000",
		2109 =>	x"0000000F",
		2110 =>	x"00000000",
		2111 =>	x"00000000",
		2112 =>	x"000F1010",
		2113 =>	x"0000000F",
		2114 =>	x"0000000F",
		2115 =>	x"10100000",
		2116 =>	x"0011110F",
		2117 =>	x"0000000F",
		2118 =>	x"00000011",
		2119 =>	x"11110000",
		2120 =>	x"000F100F",
		2121 =>	x"000F100F",
		2122 =>	x"11110011",
		2123 =>	x"10100000",
		2124 =>	x"0011110F",
		2125 =>	x"0F0F1010",
		2126 =>	x"10101111",
		2127 =>	x"11110000",
		2128 =>	x"000F100F",
		2129 =>	x"0F100F0F",
		2130 =>	x"10101011",
		2131 =>	x"10100000",
		2132 =>	x"0011110F",
		2133 =>	x"0F100F10",
		2134 =>	x"11101011",
		2135 =>	x"11110000",
		2136 =>	x"000F100F",
		2137 =>	x"0F100F10",
		2138 =>	x"11101011",
		2139 =>	x"10100000",
		2140 =>	x"0011110F",
		2141 =>	x"0F0F1011",
		2142 =>	x"11101011",
		2143 =>	x"11110000",
		2144 =>	x"000F100F",
		2145 =>	x"110F0F10",
		2146 =>	x"10101111",
		2147 =>	x"10100000",
		2148 =>	x"0011110F",
		2149 =>	x"00111111",
		2150 =>	x"11110011",
		2151 =>	x"11110000",
		2152 =>	x"000F1010",
		2153 =>	x"00000000",
		2154 =>	x"00000011",
		2155 =>	x"10100000",
		2156 =>	x"00000000",
		2157 =>	x"00000000",
		2158 =>	x"00000000",
		2159 =>	x"00000000",


--			***** MAP *****


		2160 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2161 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2162 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2163 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2164 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2165 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2166 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2167 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2168 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2169 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2170 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2171 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2172 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2173 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2174 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2175 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2176 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2177 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2178 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2179 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2180 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2181 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2182 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2183 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2184 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2185 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2186 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2187 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2188 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2189 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2190 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2191 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2192 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2193 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2194 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2195 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2196 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2197 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2198 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2199 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2200 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2201 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2202 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2203 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2204 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2205 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2206 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2207 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2208 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2209 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2210 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2211 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2212 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2213 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2214 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2215 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2216 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2217 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2218 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2219 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2220 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2221 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2222 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2223 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2224 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2225 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2226 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2227 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2228 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2229 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2230 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2231 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2232 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2233 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2234 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2235 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2236 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2237 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2238 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2239 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2240 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2241 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2242 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2243 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2244 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2245 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2246 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2247 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2248 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2249 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2250 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2251 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2252 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2253 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2254 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2255 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2256 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2257 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2258 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2259 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2260 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2261 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2262 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2263 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2264 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2265 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2266 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2267 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2268 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2269 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2270 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2271 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2272 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2273 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2274 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2275 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2276 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2277 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2278 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2279 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2280 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2281 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2282 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2283 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2284 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2285 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2286 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2287 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2288 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2289 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2290 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2291 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2292 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2293 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2294 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2295 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2296 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2297 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2298 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2299 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2300 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2301 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2302 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2303 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2304 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2305 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2306 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2307 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2308 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2309 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2310 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2311 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2312 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2313 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2314 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2315 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2316 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2317 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2318 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2319 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2320 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2321 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2322 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2323 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2324 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2325 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2326 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2327 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2328 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2329 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2330 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2331 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2332 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2333 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2334 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2335 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2336 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2337 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2338 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2339 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2340 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2341 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2342 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2343 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2344 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2345 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2346 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2347 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2348 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2349 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2350 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2351 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2352 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2353 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2354 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2355 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2356 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2357 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2358 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2359 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2360 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2361 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2362 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2363 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2364 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2365 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2366 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2367 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2368 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2369 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2370 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2371 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2372 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2373 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2374 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2375 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2376 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2377 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2378 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2379 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2380 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2381 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2382 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2383 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2384 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2385 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2386 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2387 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2388 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2389 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2390 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2391 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2392 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2393 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2394 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2395 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2396 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2397 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2398 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2399 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2400 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2401 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2402 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2403 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2404 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2405 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2406 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2407 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2408 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2409 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2410 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2411 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2412 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2413 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2414 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2415 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2416 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2417 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2418 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2419 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2420 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2421 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2422 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2423 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2424 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2425 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2426 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2427 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2428 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2429 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2430 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2431 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2432 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2433 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2434 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2435 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2436 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2437 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2438 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2439 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2440 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2441 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2442 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2443 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2444 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2445 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2446 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2447 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2448 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2449 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2450 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2451 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2452 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2453 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2454 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2455 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2456 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2457 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2458 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2459 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2460 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2461 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2462 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2463 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2464 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2465 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2466 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2467 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2468 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2469 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2470 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2471 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2472 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2473 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2474 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2475 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2476 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2477 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2478 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2479 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2480 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2481 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2482 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2483 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2484 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2485 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2486 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2487 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2488 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2489 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2490 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2491 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2492 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2493 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2494 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2495 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2496 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2497 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2498 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2499 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2500 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2501 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2502 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2503 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2504 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2505 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2506 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2507 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2508 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2509 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2510 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2511 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2512 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2513 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2514 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2515 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2516 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2517 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2518 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2519 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2520 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2521 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2522 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2523 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2524 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2525 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2526 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2527 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2528 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2529 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2530 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2531 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2532 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2533 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2534 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2535 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2536 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2537 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2538 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2539 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2540 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2541 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2542 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2543 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2544 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2545 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2546 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2547 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2548 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2549 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2550 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2551 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2552 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2553 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2554 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2555 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2556 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2557 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2558 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2559 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2560 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2561 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2562 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2563 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2564 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2565 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2566 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2567 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2568 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2569 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2570 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2571 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2572 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2573 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2574 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2575 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2576 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2577 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2578 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2579 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2580 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2581 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2582 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2583 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2584 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2585 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2586 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2587 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2588 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2589 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2590 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2591 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2592 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2593 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2594 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2595 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2596 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2597 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2598 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2599 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2600 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2601 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2602 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2603 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2604 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2605 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2606 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2607 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2608 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2609 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2610 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2611 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2612 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2613 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2614 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2615 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2616 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2617 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2618 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2619 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2620 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2621 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2622 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2623 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2624 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2625 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2626 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2627 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2628 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2629 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2630 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2631 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2632 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2633 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2634 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2635 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2636 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2637 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2638 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2639 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2640 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2641 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2642 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2643 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2644 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2645 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2646 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2647 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2648 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2649 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2650 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2651 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2652 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2653 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2654 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2655 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2656 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2657 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2658 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2659 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2660 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2661 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2662 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2663 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2664 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2665 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2666 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2667 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2668 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2669 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2670 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2671 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2672 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2673 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2674 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2675 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2676 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2677 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2678 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2679 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2680 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2681 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2682 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2683 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2684 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2685 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2686 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2687 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2688 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2689 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2690 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2691 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2692 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2693 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2694 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2695 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2696 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2697 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2698 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2699 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2700 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2701 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2702 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2703 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2704 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2705 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2706 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2707 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2708 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2709 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2710 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2711 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2712 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2713 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2714 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2715 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2716 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2717 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2718 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2719 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2720 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2721 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2722 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2723 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2724 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2725 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2726 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2727 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2728 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2729 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2730 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2731 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2732 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2733 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2734 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2735 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2736 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2737 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2738 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2739 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2740 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2741 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2742 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2743 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2744 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2745 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2746 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2747 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2748 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2749 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2750 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2751 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2752 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2753 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2754 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2755 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2756 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2757 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2758 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2759 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2760 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2761 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2762 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2763 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2764 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2765 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2766 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2767 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2768 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2769 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2770 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2771 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2772 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2773 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2774 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2775 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2776 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2777 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2778 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2779 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2780 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2781 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2782 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2783 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2784 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2785 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2786 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2787 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2788 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2789 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2790 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2791 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2792 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2793 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2794 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2795 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2796 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2797 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2798 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2799 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2800 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2801 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2802 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2803 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2804 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2805 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2806 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2807 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2808 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2809 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2810 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2811 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2812 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2813 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2814 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2815 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2816 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2817 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2818 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2819 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2820 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2821 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2822 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2823 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2824 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2825 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2826 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2827 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2828 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2829 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2830 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2831 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2832 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2833 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2834 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2835 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2836 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2837 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2838 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2839 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2840 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2841 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2842 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2843 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2844 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2845 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2846 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2847 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2848 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2849 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2850 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2851 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2852 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2853 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2854 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2855 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2856 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2857 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2858 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2859 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2860 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2861 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2862 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2863 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2864 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2865 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2866 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2867 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2868 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2869 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2870 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2871 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2872 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2873 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2874 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2875 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2876 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2877 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2878 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2879 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2880 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2881 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2882 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2883 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2884 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2885 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2886 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2887 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2888 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2889 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2890 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2891 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2892 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2893 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2894 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2895 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2896 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2897 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2898 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2899 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2900 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2901 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2902 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2903 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2904 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2905 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2906 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2907 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2908 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2909 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2910 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2911 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2912 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2913 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2914 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2915 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2916 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2917 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2918 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2919 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2920 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2921 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2922 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2923 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2924 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2925 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2926 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2927 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2928 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2929 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2930 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2931 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2932 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2933 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2934 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2935 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2936 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2937 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2938 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2939 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2940 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2941 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2942 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2943 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2944 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2945 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2946 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2947 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		2948 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2949 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2950 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2951 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2952 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2953 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2954 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2955 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2956 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2957 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2958 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2959 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2960 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2961 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2962 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2963 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2964 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2965 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2966 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2967 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		2968 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2969 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2970 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2971 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2972 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		2973 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2974 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2975 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2976 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2977 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2978 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2979 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2980 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2981 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		2982 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2983 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2984 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2985 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2986 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2987 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2988 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2989 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		2990 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		2991 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		2992 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		2993 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		2994 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2995 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2996 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2997 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2998 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2999 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3000 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3001 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3002 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3003 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3004 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3005 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3006 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3007 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3008 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3009 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3010 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3011 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3012 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3013 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3014 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3015 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3016 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3017 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3018 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3019 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3020 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3021 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3022 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3023 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3024 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3025 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3026 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3027 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3028 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3029 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3030 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3031 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3032 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3033 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3034 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3035 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3036 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3037 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3038 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3039 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3040 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3041 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3042 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3043 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3044 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3045 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3046 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3047 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3048 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3049 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3050 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3051 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3052 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3053 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3054 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3055 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3056 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3057 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3058 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3059 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3060 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3061 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3062 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3063 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3064 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3065 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3066 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3067 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3068 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3069 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3070 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3071 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3072 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3073 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3074 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3075 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3076 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3077 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3078 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3079 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3080 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3081 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3082 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3083 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3084 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3085 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3086 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3087 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3088 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3089 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3090 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3091 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3092 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3093 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3094 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3095 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3096 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3097 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3098 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3099 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3100 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3101 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3102 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3103 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3104 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3105 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3106 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3107 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3108 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3109 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3110 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3111 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3112 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3113 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3114 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3115 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3116 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3117 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3118 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3119 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3120 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3121 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3122 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3123 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3124 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3125 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3126 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3127 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3128 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3129 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3130 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3131 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3132 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3133 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3134 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3135 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3136 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3137 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3138 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3139 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3140 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3141 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3142 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3143 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3144 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3145 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3146 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3147 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3148 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3149 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3150 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3151 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3152 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3153 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3154 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3155 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3156 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3157 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3158 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3159 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3160 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3161 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3162 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3163 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3164 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3165 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3166 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3167 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3168 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3169 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3170 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3171 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3172 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3173 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3174 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3175 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3176 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3177 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3178 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3179 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3180 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3181 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3182 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3183 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3184 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3185 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3186 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3187 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3188 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3189 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3190 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3191 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3192 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3193 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3194 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3195 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3196 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3197 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3198 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3199 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3200 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3201 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3202 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3203 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3204 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3205 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3206 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3207 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3208 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3209 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3210 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3211 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3212 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3213 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3214 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3215 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3216 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3217 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3218 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3219 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3220 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3221 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3222 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3223 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3224 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3225 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3226 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3227 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3228 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3229 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3230 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3231 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3232 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3233 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3234 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3235 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3236 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3237 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3238 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3239 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3240 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3241 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3242 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3243 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3244 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3245 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3246 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3247 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3248 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3249 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3250 =>	x"000003D0", -- z: 0 rot: 0 ptr: 976
		3251 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3252 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3253 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3254 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3255 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3256 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3257 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3258 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3259 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3260 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3261 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3262 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3263 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3264 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3265 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3266 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3267 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3268 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3269 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3270 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3271 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3272 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3273 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3274 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3275 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3276 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3277 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3278 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3279 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3280 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3281 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3282 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3283 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3284 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3285 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3286 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3287 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3288 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3289 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3290 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3291 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3292 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3293 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3294 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3295 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3296 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3297 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3298 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3299 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3300 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3301 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3302 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3303 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3304 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3305 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3306 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3307 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3308 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3309 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3310 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3311 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3312 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3313 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3314 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3315 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3316 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3317 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3318 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3319 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3320 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3321 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3322 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3323 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3324 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3325 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3326 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3327 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3328 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3329 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3330 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3331 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3332 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3333 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3334 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3335 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3336 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3337 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3338 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3339 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3340 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3341 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3342 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3343 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3344 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3345 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3346 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3347 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3348 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3349 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3350 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3351 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3352 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3353 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3354 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3355 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3356 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3357 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3358 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3359 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3360 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3361 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3362 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3363 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3364 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3365 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3366 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3367 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3368 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3369 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3370 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3371 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3372 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3373 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3374 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3375 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3376 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3377 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3378 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3379 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3380 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3381 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3382 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3383 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3384 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3385 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3386 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3387 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3388 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3389 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3390 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3391 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3392 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3393 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3394 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3395 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3396 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3397 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3398 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3399 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3400 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3401 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3402 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3403 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3404 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3405 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3406 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3407 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3408 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3409 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3410 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3411 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3412 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3413 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3414 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3415 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3416 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3417 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3418 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3419 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3420 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3421 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3422 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3423 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3424 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3425 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3426 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3427 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3428 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3429 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3430 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3431 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3432 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3433 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3434 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3435 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3436 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3437 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3438 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3439 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3440 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3441 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3442 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3443 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3444 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3445 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3446 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3447 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3448 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3449 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3450 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3451 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3452 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3453 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3454 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3455 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3456 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3457 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3458 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3459 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3460 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3461 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3462 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3463 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3464 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3465 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3466 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3467 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3468 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3469 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3470 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3471 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3472 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3473 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3474 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3475 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3476 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3477 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3478 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3479 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3480 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3481 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3482 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3483 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3484 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3485 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3486 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3487 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3488 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3489 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3490 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3491 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3492 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3493 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3494 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3495 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3496 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3497 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3498 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3499 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3500 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3501 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3502 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3503 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3504 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3505 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3506 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3507 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3508 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3509 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3510 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3511 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3512 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3513 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3514 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3515 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3516 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3517 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3518 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3519 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3520 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3521 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3522 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3523 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3524 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3525 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3526 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3527 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3528 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3529 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3530 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3531 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3532 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3533 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3534 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3535 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3536 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3537 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3538 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3539 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3540 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3541 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3542 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3543 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3544 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3545 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3546 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3547 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3548 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3549 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3550 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3551 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		3552 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3553 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3554 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3555 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3556 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3557 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3558 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3559 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3560 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3561 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3562 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3563 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3564 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3565 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3566 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3567 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3568 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3569 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3570 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3571 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3572 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3573 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3574 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3575 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3576 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3577 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3578 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3579 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3580 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3581 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3582 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3583 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		3584 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3585 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3586 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3587 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3588 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3589 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3590 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3591 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3592 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3593 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3594 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3595 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3596 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3597 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3598 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3599 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3600 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3601 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3602 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3603 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3604 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3605 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3606 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3607 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3608 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3609 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3610 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3611 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3612 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3613 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3614 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3615 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3616 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3617 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3618 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3619 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3620 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3621 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3622 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3623 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3624 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3625 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3626 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3627 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3628 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3629 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3630 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3631 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3632 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3633 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3634 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3635 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3636 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3637 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3638 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3639 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3640 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3641 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3642 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3643 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3644 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3645 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3646 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3647 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3648 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3649 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3650 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3651 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3652 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3653 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3654 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3655 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3656 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3657 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3658 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3659 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3660 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3661 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3662 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3663 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3664 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3665 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3666 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3667 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3668 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3669 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3670 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3671 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3672 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3673 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3674 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3675 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3676 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3677 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3678 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3679 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3680 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3681 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3682 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3683 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3684 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3685 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3686 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3687 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3688 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3689 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3690 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3691 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3692 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3693 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3694 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3695 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3696 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3697 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3698 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3699 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3700 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3701 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3702 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3703 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3704 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3705 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3706 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3707 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3708 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3709 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3710 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3711 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3712 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3713 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3714 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3715 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3716 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3717 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3718 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3719 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3720 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3721 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3722 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3723 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3724 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3725 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3726 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3727 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3728 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3729 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3730 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3731 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3732 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3733 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3734 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3735 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3736 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3737 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3738 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3739 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3740 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3741 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3742 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3743 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3744 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3745 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3746 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3747 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3748 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3749 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3750 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3751 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3752 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3753 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3754 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3755 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3756 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3757 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3758 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3759 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3760 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3761 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3762 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3763 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3764 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3765 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3766 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3767 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3768 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3769 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3770 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3771 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3772 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3773 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3774 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3775 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3776 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3777 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3778 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3779 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3780 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3781 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3782 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3783 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3784 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3785 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3786 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3787 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3788 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3789 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3790 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3791 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3792 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3793 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3794 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3795 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3796 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3797 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3798 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3799 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3800 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3801 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3802 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3803 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3804 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3805 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3806 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3807 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3808 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3809 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3810 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3811 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3812 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3813 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3814 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3815 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3816 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3817 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3818 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3819 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3820 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3821 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3822 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3823 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3824 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3825 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3826 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3827 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3828 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3829 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3830 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3831 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3832 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3833 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3834 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3835 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3836 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3837 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3838 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3839 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3840 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3841 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3842 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3843 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3844 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3845 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3846 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3847 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3848 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3849 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3850 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3851 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3852 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3853 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3854 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3855 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3856 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3857 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3858 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3859 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3860 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3861 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3862 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3863 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3864 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3865 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3866 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3867 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3868 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3869 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3870 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3871 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3872 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3873 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3874 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3875 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3876 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3877 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3878 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3879 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3880 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3881 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3882 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3883 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3884 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3885 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3886 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3887 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3888 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3889 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3890 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3891 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3892 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3893 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3894 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3895 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3896 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3897 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3898 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3899 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3900 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3901 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3902 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3903 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3904 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3905 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3906 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3907 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3908 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3909 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3910 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3911 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3912 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3913 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3914 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3915 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3916 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3917 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3918 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3919 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3920 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3921 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3922 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3923 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3924 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3925 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3926 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3927 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3928 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3929 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3930 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3931 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3932 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3933 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3934 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3935 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3936 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3937 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3938 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3939 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3940 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3941 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3942 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3943 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3944 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3945 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3946 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3947 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3948 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3949 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3950 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3951 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3952 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3953 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3954 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3955 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3956 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3957 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3958 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3959 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3960 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3961 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3962 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3963 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3964 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3965 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3966 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3967 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3968 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3969 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3970 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3971 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3972 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3973 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3974 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3975 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3976 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3977 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3978 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3979 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3980 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3981 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3982 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3983 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		3984 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3985 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3986 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3987 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3988 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3989 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		3990 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3991 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		3992 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3993 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3994 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3995 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3996 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3997 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3998 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		3999 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4000 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4001 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4002 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4003 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4004 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4005 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4006 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4007 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4008 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4009 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4010 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4011 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4012 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4013 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4014 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4015 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4016 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4017 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4018 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4019 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4020 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4021 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4022 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4023 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4024 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4025 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4026 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4027 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4028 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4029 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4030 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4031 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4032 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4033 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4034 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4035 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4036 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4037 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4038 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4039 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4040 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4041 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4042 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4043 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4044 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4045 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4046 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4047 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4048 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4049 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4050 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4051 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4052 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4053 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4054 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4055 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4056 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4057 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4058 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4059 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4060 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4061 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4062 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4063 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4064 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4065 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4066 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4067 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4068 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4069 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4070 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4071 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4072 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4073 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4074 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4075 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4076 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4077 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4078 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4079 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4080 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4081 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4082 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4083 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4084 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4085 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4086 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4087 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4088 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4089 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4090 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4091 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4092 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4093 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4094 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4095 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4096 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4097 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4098 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4099 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4100 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4101 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4102 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4103 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4104 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4105 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4106 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4107 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4108 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4109 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4110 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4111 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4112 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4113 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4114 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4115 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4116 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4117 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4118 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4119 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4120 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4121 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4122 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4123 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4124 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4125 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4126 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4127 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4128 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4129 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4130 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4131 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4132 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4133 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4134 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4135 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4136 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4137 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4138 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4139 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4140 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4141 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4142 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4143 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4144 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4145 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4146 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4147 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4148 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4149 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4150 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4151 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4152 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4153 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4154 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4155 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4156 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4157 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4158 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4159 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4160 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4161 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4162 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4163 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4164 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4165 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4166 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4167 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4168 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4169 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4170 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4171 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4172 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4173 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4174 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4175 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4176 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4177 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4178 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4179 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4180 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4181 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4182 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4183 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4184 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4185 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4186 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4187 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4188 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4189 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4190 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4191 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4192 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4193 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4194 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4195 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4196 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4197 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4198 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4199 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4200 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4201 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4202 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4203 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4204 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4205 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4206 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4207 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4208 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4209 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4210 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4211 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4212 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4213 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4214 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4215 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4216 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4217 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4218 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4219 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4220 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4221 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4222 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4223 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4224 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4225 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4226 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4227 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4228 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4229 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4230 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4231 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4232 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4233 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4234 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4235 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4236 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4237 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4238 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4239 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4240 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4241 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4242 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4243 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4244 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4245 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4246 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4247 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4248 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4249 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4250 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4251 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4252 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4253 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4254 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4255 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4256 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4257 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4258 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4259 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4260 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4261 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4262 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4263 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4264 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4265 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4266 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4267 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4268 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4269 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4270 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4271 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4272 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4273 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4274 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4275 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4276 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4277 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4278 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4279 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4280 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4281 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4282 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4283 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4284 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4285 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4286 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4287 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4288 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4289 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4290 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4291 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4292 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4293 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4294 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4295 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4296 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4297 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4298 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4299 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4300 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4301 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4302 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4303 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4304 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4305 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4306 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4307 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4308 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4309 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4310 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4311 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4312 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4313 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4314 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4315 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4316 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4317 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4318 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4319 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4320 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4321 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4322 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4323 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4324 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4325 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4326 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4327 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4328 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4329 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4330 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4331 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4332 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4333 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4334 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4335 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4336 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4337 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4338 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4339 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4340 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4341 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4342 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4343 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4344 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4345 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4346 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4347 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4348 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4349 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4350 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4351 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4352 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4353 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4354 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4355 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4356 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4357 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4358 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4359 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4360 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4361 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4362 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4363 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4364 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4365 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4366 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4367 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4368 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4369 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4370 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4371 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4372 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4373 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4374 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4375 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4376 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4377 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4378 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4379 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4380 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4381 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4382 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4383 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4384 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4385 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4386 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4387 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4388 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4389 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4390 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4391 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4392 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4393 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4394 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4395 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4396 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4397 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4398 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4399 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4400 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4401 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4402 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4403 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4404 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4405 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4406 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4407 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4408 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4409 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4410 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4411 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4412 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4413 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4414 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4415 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4416 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4417 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4418 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4419 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4420 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4421 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4422 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4423 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4424 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4425 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4426 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4427 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4428 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4429 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4430 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4431 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4432 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4433 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4434 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4435 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4436 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4437 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4438 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4439 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4440 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4441 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4442 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4443 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4444 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4445 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4446 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4447 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4448 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4449 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4450 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4451 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4452 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4453 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4454 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4455 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4456 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4457 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4458 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4459 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4460 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4461 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4462 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4463 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4464 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4465 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4466 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4467 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4468 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4469 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4470 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4471 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4472 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4473 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4474 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4475 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4476 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4477 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4478 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4479 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4480 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4481 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4482 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4483 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4484 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4485 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4486 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4487 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4488 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4489 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4490 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4491 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4492 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4493 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4494 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4495 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4496 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4497 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4498 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4499 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4500 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4501 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4502 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4503 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4504 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4505 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4506 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4507 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4508 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4509 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4510 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4511 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4512 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4513 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4514 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4515 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4516 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4517 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4518 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4519 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4520 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		4521 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4522 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4523 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4524 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4525 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4526 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4527 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4528 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4529 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4530 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4531 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4532 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4533 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4534 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4535 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4536 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4537 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4538 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4539 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4540 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4541 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4542 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4543 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4544 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4545 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4546 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4547 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4548 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4549 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4550 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4551 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4552 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4553 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4554 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4555 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4556 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4557 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4558 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4559 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4560 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4561 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4562 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4563 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4564 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4565 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4566 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4567 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4568 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4569 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4570 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4571 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4572 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4573 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4574 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4575 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4576 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4577 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4578 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4579 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4580 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4581 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4582 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4583 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4584 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4585 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4586 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4587 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4588 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4589 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4590 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4591 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4592 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4593 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4594 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4595 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4596 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4597 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4598 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4599 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4600 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4601 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4602 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4603 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4604 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4605 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4606 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4607 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4608 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4609 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4610 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4611 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4612 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4613 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4614 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4615 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4616 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4617 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4618 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4619 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4620 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4621 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4622 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4623 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4624 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4625 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4626 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4627 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4628 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4629 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4630 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4631 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4632 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4633 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4634 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4635 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4636 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4637 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4638 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4639 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4640 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4641 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4642 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4643 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4644 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4645 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4646 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4647 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4648 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4649 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4650 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4651 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4652 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4653 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4654 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4655 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4656 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4657 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4658 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4659 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4660 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4661 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4662 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4663 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4664 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4665 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4666 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4667 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4668 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4669 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4670 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4671 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4672 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4673 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4674 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4675 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4676 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4677 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4678 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4679 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4680 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4681 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4682 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4683 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4684 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4685 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4686 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4687 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4688 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4689 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4690 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4691 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4692 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4693 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4694 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4695 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4696 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4697 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4698 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4699 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4700 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4701 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4702 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4703 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4704 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4705 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4706 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4707 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4708 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4709 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4710 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4711 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4712 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4713 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4714 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4715 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4716 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4717 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4718 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4719 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4720 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4721 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4722 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4723 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4724 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4725 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4726 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4727 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4728 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4729 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4730 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4731 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4732 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4733 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4734 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4735 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4736 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4737 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4738 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4739 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4740 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4741 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4742 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4743 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4744 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4745 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4746 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4747 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4748 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4749 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4750 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4751 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4752 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4753 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4754 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4755 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4756 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4757 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4758 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4759 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4760 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4761 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4762 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4763 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4764 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4765 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4766 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4767 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4768 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4769 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4770 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4771 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4772 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4773 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4774 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4775 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4776 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4777 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4778 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4779 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4780 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4781 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4782 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4783 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4784 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4785 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4786 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4787 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4788 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4789 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4790 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4791 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4792 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4793 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4794 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4795 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4796 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4797 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4798 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4799 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4800 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4801 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4802 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4803 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4804 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4805 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4806 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4807 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4808 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4809 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4810 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4811 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4812 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4813 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4814 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4815 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4816 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4817 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4818 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4819 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4820 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4821 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4822 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4823 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4824 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4825 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4826 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4827 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4828 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4829 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4830 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4831 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4832 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4833 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4834 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4835 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4836 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4837 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4838 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4839 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4840 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4841 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4842 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4843 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4844 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4845 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4846 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4847 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4848 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4849 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4850 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4851 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4852 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4853 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4854 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4855 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4856 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4857 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4858 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4859 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4860 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4861 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4862 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4863 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4864 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4865 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4866 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4867 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4868 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4869 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4870 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4871 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4872 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4873 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4874 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4875 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4876 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4877 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4878 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4879 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4880 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4881 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4882 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4883 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4884 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4885 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4886 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4887 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4888 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4889 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4890 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4891 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4892 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4893 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4894 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4895 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4896 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4897 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4898 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4899 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4900 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4901 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4902 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4903 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4904 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4905 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4906 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4907 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4908 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4909 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4910 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4911 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4912 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4913 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4914 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4915 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4916 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4917 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4918 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4919 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4920 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4921 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4922 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4923 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4924 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4925 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4926 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4927 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4928 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4929 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4930 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4931 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4932 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4933 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4934 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4935 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4936 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4937 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4938 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4939 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4940 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4941 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4942 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4943 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4944 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4945 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4946 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4947 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4948 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4949 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4950 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4951 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4952 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4953 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4954 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4955 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4956 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4957 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4958 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4959 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4960 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4961 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4962 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4963 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4964 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4965 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4966 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4967 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		4968 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4969 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4970 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4971 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4972 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4973 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4974 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4975 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4976 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4977 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4978 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4979 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		4980 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4981 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4982 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4983 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4984 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4985 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		4986 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4987 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		4988 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4989 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4990 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4991 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4992 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4993 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4994 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4995 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4996 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4997 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4998 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		4999 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5000 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5001 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5002 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5003 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5004 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5005 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5006 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5007 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5008 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5009 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5010 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5011 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5012 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5013 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5014 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5015 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5016 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5017 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5018 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5019 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5020 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5021 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5022 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5023 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5024 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5025 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5026 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5027 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5028 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5029 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5030 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5031 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5032 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5033 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5034 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5035 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5036 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5037 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5038 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5039 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5040 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5041 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5042 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5043 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5044 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5045 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5046 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5047 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5048 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5049 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5050 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5051 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5052 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5053 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5054 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5055 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5056 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5057 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5058 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5059 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5060 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5061 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5062 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5063 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5064 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5065 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5066 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5067 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5068 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5069 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5070 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5071 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5072 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5073 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5074 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5075 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5076 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5077 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5078 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5079 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5080 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5081 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5082 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5083 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5084 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5085 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5086 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5087 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5088 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5089 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5090 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5091 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5092 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5093 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5094 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5095 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5096 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5097 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5098 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5099 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5100 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5101 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5102 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5103 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5104 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5105 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5106 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5107 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5108 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5109 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5110 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5111 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5112 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5113 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5114 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5115 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5116 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5117 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5118 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5119 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5120 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5121 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5122 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5123 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5124 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5125 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5126 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5127 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5128 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5129 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5130 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5131 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5132 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5133 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5134 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5135 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5136 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5137 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5138 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5139 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5140 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5141 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5142 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5143 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5144 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5145 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5146 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5147 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5148 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5149 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5150 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5151 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5152 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5153 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5154 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5155 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5156 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5157 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5158 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5159 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5160 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5161 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5162 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5163 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5164 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5165 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5166 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5167 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5168 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5169 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5170 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5171 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5172 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5173 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5174 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5175 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5176 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5177 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5178 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5179 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5180 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5181 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5182 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5183 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5184 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5185 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5186 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5187 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5188 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5189 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5190 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5191 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5192 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5193 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5194 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5195 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5196 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5197 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5198 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5199 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5200 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5201 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5202 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5203 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5204 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5205 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5206 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5207 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5208 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5209 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5210 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5211 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5212 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5213 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5214 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5215 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5216 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5217 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5218 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5219 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5220 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5221 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5222 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5223 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5224 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5225 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5226 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5227 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5228 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5229 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5230 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5231 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5232 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5233 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5234 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5235 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5236 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5237 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5238 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5239 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5240 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5241 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5242 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5243 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5244 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5245 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5246 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5247 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5248 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5249 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5250 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5251 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5252 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5253 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5254 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5255 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5256 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5257 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5258 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5259 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5260 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5261 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5262 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5263 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5264 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5265 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5266 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5267 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5268 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5269 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5270 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5271 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5272 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5273 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5274 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5275 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5276 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5277 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5278 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5279 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5280 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5281 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5282 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5283 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5284 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5285 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5286 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5287 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5288 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5289 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5290 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5291 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5292 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5293 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5294 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5295 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5296 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5297 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5298 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5299 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5300 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5301 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5302 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5303 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5304 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5305 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5306 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5307 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5308 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5309 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5310 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5311 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5312 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5313 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5314 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5315 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5316 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5317 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5318 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5319 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5320 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5321 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5322 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5323 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5324 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5325 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5326 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5327 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5328 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5329 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5330 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5331 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5332 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5333 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5334 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5335 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5336 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5337 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5338 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5339 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5340 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5341 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5342 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5343 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5344 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5345 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5346 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5347 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5348 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5349 =>	x"00000420", -- z: 0 rot: 0 ptr: 1056
		5350 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5351 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5352 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5353 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5354 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5355 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5356 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5357 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5358 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5359 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5360 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5361 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5362 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5363 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5364 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5365 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5366 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5367 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5368 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5369 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5370 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5371 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5372 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5373 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5374 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5375 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5376 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5377 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5378 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5379 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5380 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5381 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5382 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5383 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5384 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5385 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5386 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5387 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5388 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5389 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5390 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5391 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5392 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5393 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5394 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5395 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5396 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5397 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5398 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5399 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5400 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5401 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5402 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5403 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5404 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5405 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5406 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5407 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5408 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5409 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5410 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5411 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5412 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5413 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5414 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5415 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5416 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5417 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5418 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5419 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5420 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5421 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5422 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5423 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5424 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5425 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5426 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5427 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5428 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5429 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5430 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5431 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5432 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5433 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5434 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5435 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5436 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5437 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5438 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5439 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5440 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5441 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5442 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5443 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5444 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5445 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5446 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5447 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5448 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5449 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5450 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5451 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5452 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5453 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5454 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5455 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5456 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5457 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5458 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5459 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5460 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5461 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5462 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5463 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5464 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5465 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5466 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5467 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5468 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5469 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5470 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5471 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5472 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5473 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5474 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5475 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5476 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5477 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5478 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5479 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5480 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5481 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5482 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5483 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5484 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5485 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5486 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5487 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5488 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5489 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5490 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5491 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5492 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5493 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5494 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5495 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5496 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5497 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5498 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5499 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5500 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5501 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5502 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5503 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5504 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5505 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5506 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5507 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5508 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5509 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5510 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5511 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5512 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5513 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5514 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5515 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5516 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5517 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5518 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5519 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5520 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5521 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5522 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5523 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5524 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5525 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5526 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5527 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5528 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5529 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5530 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5531 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5532 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5533 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5534 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5535 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5536 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5537 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5538 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5539 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5540 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5541 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5542 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5543 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5544 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5545 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5546 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5547 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5548 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5549 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5550 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5551 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5552 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5553 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5554 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5555 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5556 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5557 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5558 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5559 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5560 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5561 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5562 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5563 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5564 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5565 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5566 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5567 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5568 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5569 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5570 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5571 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5572 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5573 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5574 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5575 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5576 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5577 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5578 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5579 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5580 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5581 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5582 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5583 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5584 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5585 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5586 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5587 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5588 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5589 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5590 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5591 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5592 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5593 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5594 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5595 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5596 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5597 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5598 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5599 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5600 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5601 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5602 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5603 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5604 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5605 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5606 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5607 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5608 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5609 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5610 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5611 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5612 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5613 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5614 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5615 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5616 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5617 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5618 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5619 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5620 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5621 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5622 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5623 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5624 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5625 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5626 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5627 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5628 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5629 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5630 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5631 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5632 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5633 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5634 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5635 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5636 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5637 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5638 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5639 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5640 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5641 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5642 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5643 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5644 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5645 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5646 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5647 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5648 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5649 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5650 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5651 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5652 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5653 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5654 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5655 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5656 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5657 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5658 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5659 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5660 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5661 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5662 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5663 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5664 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5665 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5666 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5667 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5668 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5669 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5670 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5671 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5672 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5673 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5674 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5675 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5676 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5677 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5678 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5679 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5680 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5681 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5682 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5683 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5684 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5685 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5686 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5687 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5688 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5689 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5690 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5691 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5692 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5693 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5694 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5695 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5696 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5697 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5698 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5699 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5700 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5701 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5702 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5703 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5704 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5705 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5706 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5707 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5708 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5709 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5710 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5711 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5712 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5713 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5714 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5715 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5716 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5717 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5718 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5719 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5720 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5721 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		5722 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5723 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5724 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5725 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5726 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5727 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5728 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5729 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5730 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5731 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5732 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5733 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5734 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5735 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5736 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5737 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5738 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5739 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5740 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5741 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5742 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5743 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5744 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5745 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5746 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5747 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5748 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5749 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5750 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5751 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5752 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5753 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5754 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5755 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5756 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5757 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5758 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5759 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5760 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5761 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5762 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5763 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5764 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5765 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5766 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5767 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5768 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5769 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5770 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5771 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5772 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5773 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5774 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5775 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5776 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5777 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5778 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5779 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5780 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5781 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5782 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5783 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5784 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5785 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5786 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5787 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5788 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5789 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5790 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5791 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5792 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5793 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5794 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5795 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5796 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5797 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5798 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5799 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5800 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5801 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5802 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5803 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5804 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5805 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5806 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5807 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5808 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5809 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5810 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5811 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5812 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5813 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5814 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5815 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5816 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5817 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5818 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5819 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5820 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5821 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5822 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5823 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5824 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5825 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5826 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5827 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5828 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5829 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5830 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5831 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5832 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5833 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5834 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5835 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5836 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5837 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5838 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5839 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5840 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5841 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5842 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5843 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5844 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5845 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5846 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5847 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5848 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5849 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5850 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5851 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5852 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5853 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5854 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5855 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5856 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5857 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5858 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5859 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5860 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5861 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5862 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5863 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5864 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5865 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5866 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5867 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5868 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5869 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5870 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5871 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5872 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5873 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5874 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5875 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5876 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5877 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5878 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5879 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5880 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5881 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5882 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5883 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5884 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5885 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5886 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5887 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5888 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5889 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5890 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5891 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5892 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5893 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5894 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5895 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5896 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5897 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5898 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5899 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5900 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5901 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5902 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5903 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5904 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5905 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5906 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5907 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5908 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5909 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5910 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5911 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5912 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5913 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5914 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5915 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5916 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5917 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5918 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5919 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5920 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5921 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5922 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5923 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5924 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5925 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5926 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5927 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5928 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5929 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5930 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5931 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5932 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5933 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5934 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5935 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5936 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5937 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5938 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5939 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5940 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5941 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5942 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5943 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5944 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5945 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5946 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5947 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5948 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5949 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5950 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5951 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5952 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5953 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5954 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5955 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5956 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5957 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5958 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5959 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5960 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5961 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5962 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5963 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5964 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5965 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5966 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5967 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5968 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5969 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5970 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5971 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5972 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5973 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5974 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5975 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5976 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5977 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5978 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5979 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5980 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5981 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5982 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5983 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5984 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5985 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		5986 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5987 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		5988 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5989 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5990 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5991 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		5992 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5993 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5994 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5995 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5996 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5997 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5998 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		5999 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6000 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6001 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6002 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6003 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6004 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6005 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6006 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6007 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6008 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6009 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6010 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6011 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6012 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6013 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6014 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6015 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6016 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6017 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6018 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6019 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6020 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6021 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6022 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6023 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6024 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6025 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6026 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6027 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6028 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6029 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6030 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6031 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6032 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6033 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6034 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6035 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6036 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6037 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6038 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6039 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6040 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6041 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6042 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6043 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6044 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6045 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6046 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6047 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6048 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6049 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6050 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6051 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6052 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6053 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6054 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6055 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6056 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6057 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6058 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6059 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6060 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6061 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6062 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6063 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6064 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6065 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6066 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6067 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6068 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6069 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6070 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6071 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6072 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6073 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6074 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6075 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6076 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6077 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6078 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6079 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6080 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6081 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6082 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6083 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6084 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6085 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6086 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6087 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6088 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6089 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6090 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6091 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6092 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6093 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6094 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6095 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6096 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6097 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6098 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6099 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6100 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6101 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6102 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6103 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6104 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6105 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6106 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6107 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6108 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6109 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6110 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6111 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6112 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6113 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6114 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6115 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6116 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6117 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6118 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6119 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6120 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6121 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6122 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6123 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6124 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6125 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6126 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6127 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6128 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6129 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6130 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6131 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6132 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6133 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6134 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6135 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6136 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6137 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6138 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6139 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6140 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6141 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6142 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6143 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6144 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6145 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6146 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6147 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6148 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6149 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6150 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6151 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6152 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6153 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6154 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6155 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6156 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6157 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6158 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6159 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6160 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6161 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6162 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6163 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6164 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6165 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6166 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6167 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6168 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6169 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6170 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6171 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6172 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6173 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6174 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6175 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6176 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6177 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6178 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6179 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6180 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6181 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6182 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6183 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6184 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6185 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6186 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6187 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6188 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6189 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6190 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6191 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6192 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6193 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6194 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6195 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6196 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6197 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6198 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6199 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6200 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6201 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6202 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6203 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6204 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6205 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6206 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6207 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6208 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6209 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6210 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6211 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6212 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6213 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6214 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6215 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6216 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6217 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6218 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6219 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6220 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6221 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6222 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6223 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6224 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6225 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6226 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6227 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6228 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6229 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6230 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6231 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6232 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6233 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6234 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6235 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6236 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6237 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6238 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6239 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6240 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6241 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6242 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6243 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6244 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6245 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6246 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6247 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6248 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6249 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6250 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6251 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6252 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6253 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6254 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6255 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6256 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6257 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6258 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6259 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6260 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6261 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6262 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6263 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6264 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6265 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6266 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6267 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6268 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6269 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6270 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6271 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6272 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6273 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6274 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6275 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6276 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6277 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6278 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6279 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6280 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6281 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6282 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6283 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6284 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6285 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6286 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6287 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6288 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6289 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6290 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6291 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6292 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6293 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6294 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6295 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6296 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6297 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6298 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6299 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6300 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6301 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6302 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6303 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6304 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6305 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6306 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6307 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6308 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6309 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6310 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6311 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6312 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6313 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6314 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6315 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6316 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6317 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6318 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6319 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6320 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6321 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6322 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6323 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6324 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6325 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6326 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6327 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6328 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6329 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6330 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6331 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6332 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6333 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6334 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6335 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6336 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6337 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6338 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6339 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6340 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6341 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6342 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6343 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6344 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6345 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6346 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6347 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6348 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6349 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6350 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6351 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6352 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6353 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6354 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6355 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6356 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6357 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6358 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6359 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6360 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6361 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6362 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6363 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6364 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6365 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6366 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6367 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6368 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6369 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6370 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6371 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6372 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6373 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6374 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6375 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6376 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6377 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6378 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6379 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6380 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6381 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6382 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6383 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6384 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6385 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6386 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6387 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6388 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6389 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6390 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6391 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6392 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6393 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6394 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6395 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6396 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6397 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6398 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6399 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6400 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6401 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6402 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6403 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6404 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6405 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6406 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6407 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6408 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6409 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6410 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6411 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6412 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6413 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6414 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6415 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6416 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6417 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6418 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6419 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6420 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6421 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6422 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6423 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6424 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6425 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6426 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6427 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6428 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6429 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6430 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6431 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6432 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6433 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6434 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6435 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6436 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6437 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6438 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6439 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6440 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6441 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6442 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6443 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6444 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6445 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6446 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6447 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6448 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6449 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6450 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6451 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6452 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6453 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6454 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6455 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6456 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6457 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6458 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6459 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6460 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6461 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6462 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6463 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6464 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6465 =>	x"010003E0", -- z: 1 rot: 0 ptr: 992
		6466 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6467 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6468 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6469 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6470 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6471 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6472 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6473 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6474 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6475 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6476 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6477 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6478 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6479 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6480 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6481 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6482 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6483 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6484 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6485 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6486 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6487 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6488 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6489 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6490 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6491 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6492 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6493 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6494 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6495 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6496 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6497 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6498 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6499 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6500 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6501 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6502 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6503 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6504 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6505 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6506 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6507 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6508 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6509 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6510 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6511 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6512 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6513 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6514 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6515 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6516 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6517 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6518 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6519 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6520 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6521 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6522 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6523 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6524 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6525 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6526 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6527 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6528 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6529 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6530 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6531 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6532 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6533 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6534 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6535 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6536 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6537 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6538 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6539 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6540 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6541 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6542 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6543 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6544 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6545 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6546 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6547 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6548 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6549 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6550 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6551 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6552 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6553 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6554 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6555 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6556 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6557 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6558 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6559 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6560 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6561 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6562 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6563 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6564 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6565 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6566 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6567 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6568 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6569 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6570 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6571 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6572 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6573 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6574 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6575 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6576 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6577 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6578 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6579 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6580 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6581 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6582 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6583 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6584 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6585 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6586 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6587 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6588 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6589 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6590 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6591 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6592 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6593 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6594 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6595 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6596 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6597 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6598 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6599 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6600 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6601 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6602 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6603 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6604 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6605 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6606 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6607 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6608 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6609 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6610 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6611 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6612 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6613 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6614 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6615 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6616 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6617 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6618 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6619 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6620 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6621 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6622 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6623 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6624 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6625 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6626 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6627 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6628 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6629 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6630 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6631 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6632 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6633 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6634 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6635 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6636 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6637 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6638 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6639 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6640 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6641 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6642 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6643 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6644 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6645 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6646 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6647 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6648 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6649 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6650 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6651 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6652 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6653 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6654 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6655 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6656 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6657 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6658 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6659 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6660 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6661 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6662 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6663 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6664 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6665 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6666 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6667 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6668 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6669 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6670 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6671 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6672 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6673 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6674 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6675 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6676 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6677 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6678 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6679 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6680 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6681 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6682 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6683 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6684 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6685 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6686 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6687 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6688 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6689 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6690 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6691 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6692 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6693 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6694 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6695 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6696 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6697 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6698 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6699 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6700 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6701 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6702 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6703 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6704 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6705 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6706 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6707 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6708 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6709 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6710 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6711 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6712 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6713 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6714 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6715 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6716 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6717 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6718 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6719 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6720 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6721 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6722 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6723 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6724 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6725 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6726 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6727 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6728 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6729 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6730 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6731 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6732 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6733 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6734 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6735 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6736 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6737 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6738 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6739 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6740 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6741 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6742 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6743 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6744 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6745 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6746 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6747 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6748 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6749 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6750 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6751 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6752 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6753 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6754 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6755 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6756 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6757 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6758 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6759 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6760 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6761 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6762 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6763 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6764 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6765 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6766 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6767 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6768 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6769 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6770 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6771 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6772 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6773 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6774 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6775 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6776 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6777 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6778 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6779 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6780 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6781 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6782 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6783 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6784 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6785 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6786 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6787 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6788 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6789 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6790 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6791 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6792 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6793 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6794 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6795 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6796 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6797 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6798 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6799 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6800 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6801 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6802 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6803 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6804 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6805 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6806 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6807 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6808 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6809 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6810 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6811 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6812 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6813 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6814 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6815 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6816 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6817 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6818 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6819 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6820 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6821 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6822 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6823 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6824 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6825 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6826 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6827 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6828 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6829 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6830 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6831 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6832 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6833 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6834 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6835 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6836 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6837 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6838 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6839 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6840 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6841 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6842 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6843 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6844 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6845 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6846 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6847 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6848 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6849 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6850 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6851 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6852 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6853 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6854 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6855 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6856 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6857 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6858 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6859 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6860 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6861 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6862 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6863 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6864 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6865 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6866 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6867 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6868 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6869 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6870 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6871 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6872 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6873 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6874 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6875 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6876 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6877 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6878 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6879 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6880 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6881 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6882 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6883 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6884 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6885 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6886 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6887 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6888 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6889 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6890 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6891 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6892 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6893 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6894 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6895 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6896 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6897 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6898 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6899 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6900 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6901 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6902 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6903 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6904 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6905 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6906 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6907 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6908 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6909 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6910 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6911 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6912 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6913 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6914 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6915 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6916 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6917 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6918 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6919 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6920 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6921 =>	x"010003B0", -- z: 1 rot: 0 ptr: 944
		6922 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6923 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6924 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6925 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6926 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6927 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6928 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6929 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6930 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6931 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6932 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6933 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6934 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6935 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6936 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6937 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6938 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6939 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6940 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6941 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6942 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6943 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6944 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6945 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6946 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6947 =>	x"020003C0", -- z: 2 rot: 0 ptr: 960
		6948 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6949 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6950 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6951 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		6952 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6953 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6954 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6955 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6956 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6957 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6958 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		6959 =>	x"000003A0", -- z: 0 rot: 0 ptr: 928
		others => x"00000000"
	);

begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;