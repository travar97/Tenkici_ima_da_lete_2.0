
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);
	
	port
	(
		clk_i    : in  	std_logic;
		addr_i	: in  	std_logic_vector( ADDR_WIDTH-1 downto 0 );
		data_o	: out	std_logic_vector( DATA_WIDTH-1 downto 0 )
	);
end entity ram;

architecture arch of ram is

	type	ram_t is array ( 0 to 2**ADDR_WIDTH-1 ) of std_logic_vector( DATA_WIDTH-1 downto 0 );
	
-- GENERATED BY BC_MEM_PACKER
-- DATE: Tue Jun 02 15:48:57 2015

	signal mem : ram_t := (


--			***** COLOR PALLETE *****


		0 =>	"10000000000000000000000000000000", -- R: 128 G: 0 B: 0
		1 =>	"01100000011000001000000000000000", -- R: 96 G: 96 B: 128
		2 =>	"10100000010000000000000000000000", -- R: 160 G: 64 B: 0
		3 =>	"00000000000000000000000000000000", -- R: 0 G: 0 B: 0
		4 =>	"10100000101000001010010000000000", -- R: 160 G: 160 B: 164
		5 =>	"00000000011000000000000000000000", -- R: 0 G: 96 B: 0
		6 =>	"00000000010000000000000000000000", -- R: 0 G: 64 B: 0
		7 =>	"10000000111000000000000000000000", -- R: 128 G: 224 B: 0
		8 =>	"11111111111111111111111100000000", -- R: 255 G: 255 B: 255
		9 =>	"11000011110000111100001100000000", -- R: 195 G: 195 B: 195
		10 =>	"11000100110001001100010000000000", -- R: 196 G: 196 B: 196
		11 =>	"11000010110000101100001000000000", -- R: 194 G: 194 B: 194
		12 =>	"01000000010000001100000000000000", -- R: 64 G: 64 B: 192
		13 =>	"10100110110010101111000000000000", -- R: 166 G: 202 B: 240
		14 =>	"00000000010000000100000000000000", -- R: 0 G: 64 B: 64
		15 =>	"01100000000000001000000000000000", -- R: 96 G: 0 B: 128
		16 =>	"11000000010000000100000000000000", -- R: 192 G: 64 B: 64
		17 =>	"11100000111000001000000000000000", -- R: 224 G: 224 B: 128
		18 =>	"11100000101000000100000000000000", -- R: 224 G: 160 B: 64
		19 =>	"01100000011000000000000000000000", -- R: 96 G: 96 B: 0
		20 =>	"00000000000000000000000000000000", -- Unused
		21 =>	"00000000000000000000000000000000", -- Unused
		22 =>	"00000000000000000000000000000000", -- Unused
		23 =>	"00000000000000000000000000000000", -- Unused
		24 =>	"00000000000000000000000000000000", -- Unused
		25 =>	"00000000000000000000000000000000", -- Unused
		26 =>	"00000000000000000000000000000000", -- Unused
		27 =>	"00000000000000000000000000000000", -- Unused
		28 =>	"00000000000000000000000000000000", -- Unused
		29 =>	"00000000000000000000000000000000", -- Unused
		30 =>	"00000000000000000000000000000000", -- Unused
		31 =>	"00000000000000000000000000000000", -- Unused
		32 =>	"00000000000000000000000000000000", -- Unused
		33 =>	"00000000000000000000000000000000", -- Unused
		34 =>	"00000000000000000000000000000000", -- Unused
		35 =>	"00000000000000000000000000000000", -- Unused
		36 =>	"00000000000000000000000000000000", -- Unused
		37 =>	"00000000000000000000000000000000", -- Unused
		38 =>	"00000000000000000000000000000000", -- Unused
		39 =>	"00000000000000000000000000000000", -- Unused
		40 =>	"00000000000000000000000000000000", -- Unused
		41 =>	"00000000000000000000000000000000", -- Unused
		42 =>	"00000000000000000000000000000000", -- Unused
		43 =>	"00000000000000000000000000000000", -- Unused
		44 =>	"00000000000000000000000000000000", -- Unused
		45 =>	"00000000000000000000000000000000", -- Unused
		46 =>	"00000000000000000000000000000000", -- Unused
		47 =>	"00000000000000000000000000000000", -- Unused
		48 =>	"00000000000000000000000000000000", -- Unused
		49 =>	"00000000000000000000000000000000", -- Unused
		50 =>	"00000000000000000000000000000000", -- Unused
		51 =>	"00000000000000000000000000000000", -- Unused
		52 =>	"00000000000000000000000000000000", -- Unused
		53 =>	"00000000000000000000000000000000", -- Unused
		54 =>	"00000000000000000000000000000000", -- Unused
		55 =>	"00000000000000000000000000000000", -- Unused
		56 =>	"00000000000000000000000000000000", -- Unused
		57 =>	"00000000000000000000000000000000", -- Unused
		58 =>	"00000000000000000000000000000000", -- Unused
		59 =>	"00000000000000000000000000000000", -- Unused
		60 =>	"00000000000000000000000000000000", -- Unused
		61 =>	"00000000000000000000000000000000", -- Unused
		62 =>	"00000000000000000000000000000000", -- Unused
		63 =>	"00000000000000000000000000000000", -- Unused
		64 =>	"00000000000000000000000000000000", -- Unused
		65 =>	"00000000000000000000000000000000", -- Unused
		66 =>	"00000000000000000000000000000000", -- Unused
		67 =>	"00000000000000000000000000000000", -- Unused
		68 =>	"00000000000000000000000000000000", -- Unused
		69 =>	"00000000000000000000000000000000", -- Unused
		70 =>	"00000000000000000000000000000000", -- Unused
		71 =>	"00000000000000000000000000000000", -- Unused
		72 =>	"00000000000000000000000000000000", -- Unused
		73 =>	"00000000000000000000000000000000", -- Unused
		74 =>	"00000000000000000000000000000000", -- Unused
		75 =>	"00000000000000000000000000000000", -- Unused
		76 =>	"00000000000000000000000000000000", -- Unused
		77 =>	"00000000000000000000000000000000", -- Unused
		78 =>	"00000000000000000000000000000000", -- Unused
		79 =>	"00000000000000000000000000000000", -- Unused
		80 =>	"00000000000000000000000000000000", -- Unused
		81 =>	"00000000000000000000000000000000", -- Unused
		82 =>	"00000000000000000000000000000000", -- Unused
		83 =>	"00000000000000000000000000000000", -- Unused
		84 =>	"00000000000000000000000000000000", -- Unused
		85 =>	"00000000000000000000000000000000", -- Unused
		86 =>	"00000000000000000000000000000000", -- Unused
		87 =>	"00000000000000000000000000000000", -- Unused
		88 =>	"00000000000000000000000000000000", -- Unused
		89 =>	"00000000000000000000000000000000", -- Unused
		90 =>	"00000000000000000000000000000000", -- Unused
		91 =>	"00000000000000000000000000000000", -- Unused
		92 =>	"00000000000000000000000000000000", -- Unused
		93 =>	"00000000000000000000000000000000", -- Unused
		94 =>	"00000000000000000000000000000000", -- Unused
		95 =>	"00000000000000000000000000000000", -- Unused
		96 =>	"00000000000000000000000000000000", -- Unused
		97 =>	"00000000000000000000000000000000", -- Unused
		98 =>	"00000000000000000000000000000000", -- Unused
		99 =>	"00000000000000000000000000000000", -- Unused
		100 =>	"00000000000000000000000000000000", -- Unused
		101 =>	"00000000000000000000000000000000", -- Unused
		102 =>	"00000000000000000000000000000000", -- Unused
		103 =>	"00000000000000000000000000000000", -- Unused
		104 =>	"00000000000000000000000000000000", -- Unused
		105 =>	"00000000000000000000000000000000", -- Unused
		106 =>	"00000000000000000000000000000000", -- Unused
		107 =>	"00000000000000000000000000000000", -- Unused
		108 =>	"00000000000000000000000000000000", -- Unused
		109 =>	"00000000000000000000000000000000", -- Unused
		110 =>	"00000000000000000000000000000000", -- Unused
		111 =>	"00000000000000000000000000000000", -- Unused
		112 =>	"00000000000000000000000000000000", -- Unused
		113 =>	"00000000000000000000000000000000", -- Unused
		114 =>	"00000000000000000000000000000000", -- Unused
		115 =>	"00000000000000000000000000000000", -- Unused
		116 =>	"00000000000000000000000000000000", -- Unused
		117 =>	"00000000000000000000000000000000", -- Unused
		118 =>	"00000000000000000000000000000000", -- Unused
		119 =>	"00000000000000000000000000000000", -- Unused
		120 =>	"00000000000000000000000000000000", -- Unused
		121 =>	"00000000000000000000000000000000", -- Unused
		122 =>	"00000000000000000000000000000000", -- Unused
		123 =>	"00000000000000000000000000000000", -- Unused
		124 =>	"00000000000000000000000000000000", -- Unused
		125 =>	"00000000000000000000000000000000", -- Unused
		126 =>	"00000000000000000000000000000000", -- Unused
		127 =>	"00000000000000000000000000000000", -- Unused
		128 =>	"00000000000000000000000000000000", -- Unused
		129 =>	"00000000000000000000000000000000", -- Unused
		130 =>	"00000000000000000000000000000000", -- Unused
		131 =>	"00000000000000000000000000000000", -- Unused
		132 =>	"00000000000000000000000000000000", -- Unused
		133 =>	"00000000000000000000000000000000", -- Unused
		134 =>	"00000000000000000000000000000000", -- Unused
		135 =>	"00000000000000000000000000000000", -- Unused
		136 =>	"00000000000000000000000000000000", -- Unused
		137 =>	"00000000000000000000000000000000", -- Unused
		138 =>	"00000000000000000000000000000000", -- Unused
		139 =>	"00000000000000000000000000000000", -- Unused
		140 =>	"00000000000000000000000000000000", -- Unused
		141 =>	"00000000000000000000000000000000", -- Unused
		142 =>	"00000000000000000000000000000000", -- Unused
		143 =>	"00000000000000000000000000000000", -- Unused
		144 =>	"00000000000000000000000000000000", -- Unused
		145 =>	"00000000000000000000000000000000", -- Unused
		146 =>	"00000000000000000000000000000000", -- Unused
		147 =>	"00000000000000000000000000000000", -- Unused
		148 =>	"00000000000000000000000000000000", -- Unused
		149 =>	"00000000000000000000000000000000", -- Unused
		150 =>	"00000000000000000000000000000000", -- Unused
		151 =>	"00000000000000000000000000000000", -- Unused
		152 =>	"00000000000000000000000000000000", -- Unused
		153 =>	"00000000000000000000000000000000", -- Unused
		154 =>	"00000000000000000000000000000000", -- Unused
		155 =>	"00000000000000000000000000000000", -- Unused
		156 =>	"00000000000000000000000000000000", -- Unused
		157 =>	"00000000000000000000000000000000", -- Unused
		158 =>	"00000000000000000000000000000000", -- Unused
		159 =>	"00000000000000000000000000000000", -- Unused
		160 =>	"00000000000000000000000000000000", -- Unused
		161 =>	"00000000000000000000000000000000", -- Unused
		162 =>	"00000000000000000000000000000000", -- Unused
		163 =>	"00000000000000000000000000000000", -- Unused
		164 =>	"00000000000000000000000000000000", -- Unused
		165 =>	"00000000000000000000000000000000", -- Unused
		166 =>	"00000000000000000000000000000000", -- Unused
		167 =>	"00000000000000000000000000000000", -- Unused
		168 =>	"00000000000000000000000000000000", -- Unused
		169 =>	"00000000000000000000000000000000", -- Unused
		170 =>	"00000000000000000000000000000000", -- Unused
		171 =>	"00000000000000000000000000000000", -- Unused
		172 =>	"00000000000000000000000000000000", -- Unused
		173 =>	"00000000000000000000000000000000", -- Unused
		174 =>	"00000000000000000000000000000000", -- Unused
		175 =>	"00000000000000000000000000000000", -- Unused
		176 =>	"00000000000000000000000000000000", -- Unused
		177 =>	"00000000000000000000000000000000", -- Unused
		178 =>	"00000000000000000000000000000000", -- Unused
		179 =>	"00000000000000000000000000000000", -- Unused
		180 =>	"00000000000000000000000000000000", -- Unused
		181 =>	"00000000000000000000000000000000", -- Unused
		182 =>	"00000000000000000000000000000000", -- Unused
		183 =>	"00000000000000000000000000000000", -- Unused
		184 =>	"00000000000000000000000000000000", -- Unused
		185 =>	"00000000000000000000000000000000", -- Unused
		186 =>	"00000000000000000000000000000000", -- Unused
		187 =>	"00000000000000000000000000000000", -- Unused
		188 =>	"00000000000000000000000000000000", -- Unused
		189 =>	"00000000000000000000000000000000", -- Unused
		190 =>	"00000000000000000000000000000000", -- Unused
		191 =>	"00000000000000000000000000000000", -- Unused
		192 =>	"00000000000000000000000000000000", -- Unused
		193 =>	"00000000000000000000000000000000", -- Unused
		194 =>	"00000000000000000000000000000000", -- Unused
		195 =>	"00000000000000000000000000000000", -- Unused
		196 =>	"00000000000000000000000000000000", -- Unused
		197 =>	"00000000000000000000000000000000", -- Unused
		198 =>	"00000000000000000000000000000000", -- Unused
		199 =>	"00000000000000000000000000000000", -- Unused
		200 =>	"00000000000000000000000000000000", -- Unused
		201 =>	"00000000000000000000000000000000", -- Unused
		202 =>	"00000000000000000000000000000000", -- Unused
		203 =>	"00000000000000000000000000000000", -- Unused
		204 =>	"00000000000000000000000000000000", -- Unused
		205 =>	"00000000000000000000000000000000", -- Unused
		206 =>	"00000000000000000000000000000000", -- Unused
		207 =>	"00000000000000000000000000000000", -- Unused
		208 =>	"00000000000000000000000000000000", -- Unused
		209 =>	"00000000000000000000000000000000", -- Unused
		210 =>	"00000000000000000000000000000000", -- Unused
		211 =>	"00000000000000000000000000000000", -- Unused
		212 =>	"00000000000000000000000000000000", -- Unused
		213 =>	"00000000000000000000000000000000", -- Unused
		214 =>	"00000000000000000000000000000000", -- Unused
		215 =>	"00000000000000000000000000000000", -- Unused
		216 =>	"00000000000000000000000000000000", -- Unused
		217 =>	"00000000000000000000000000000000", -- Unused
		218 =>	"00000000000000000000000000000000", -- Unused
		219 =>	"00000000000000000000000000000000", -- Unused
		220 =>	"00000000000000000000000000000000", -- Unused
		221 =>	"00000000000000000000000000000000", -- Unused
		222 =>	"00000000000000000000000000000000", -- Unused
		223 =>	"00000000000000000000000000000000", -- Unused
		224 =>	"00000000000000000000000000000000", -- Unused
		225 =>	"00000000000000000000000000000000", -- Unused
		226 =>	"00000000000000000000000000000000", -- Unused
		227 =>	"00000000000000000000000000000000", -- Unused
		228 =>	"00000000000000000000000000000000", -- Unused
		229 =>	"00000000000000000000000000000000", -- Unused
		230 =>	"00000000000000000000000000000000", -- Unused
		231 =>	"00000000000000000000000000000000", -- Unused
		232 =>	"00000000000000000000000000000000", -- Unused
		233 =>	"00000000000000000000000000000000", -- Unused
		234 =>	"00000000000000000000000000000000", -- Unused
		235 =>	"00000000000000000000000000000000", -- Unused
		236 =>	"00000000000000000000000000000000", -- Unused
		237 =>	"00000000000000000000000000000000", -- Unused
		238 =>	"00000000000000000000000000000000", -- Unused
		239 =>	"00000000000000000000000000000000", -- Unused
		240 =>	"00000000000000000000000000000000", -- Unused
		241 =>	"00000000000000000000000000000000", -- Unused
		242 =>	"00000000000000000000000000000000", -- Unused
		243 =>	"00000000000000000000000000000000", -- Unused
		244 =>	"00000000000000000000000000000000", -- Unused
		245 =>	"00000000000000000000000000000000", -- Unused
		246 =>	"00000000000000000000000000000000", -- Unused
		247 =>	"00000000000000000000000000000000", -- Unused
		248 =>	"00000000000000000000000000000000", -- Unused
		249 =>	"00000000000000000000000000000000", -- Unused
		250 =>	"00000000000000000000000000000000", -- Unused
		251 =>	"00000000000000000000000000000000", -- Unused
		252 =>	"00000000000000000000000000000000", -- Unused
		253 =>	"00000000000000000000000000000000", -- Unused
		254 =>	"00000000000000000000000000000000", -- Unused
		255 =>	"00000000000000000000000000000000", -- Unused


--			***** 8x8 IMAGES *****


		256 =>	"00000000000000000000000000000000", -- IMG_8x8_BRICK
		257 =>	"00000001000000000000000000000000",
		258 =>	"00000010000000100000001000000010",
		259 =>	"00000001000000000000001000000010",
		260 =>	"00000010000000100000001000000010",
		261 =>	"00000001000000000000001000000010",
		262 =>	"00000001000000010000000100000001",
		263 =>	"00000001000000010000000100000001",
		264 =>	"00000001000000000000000000000000",
		265 =>	"00000000000000000000000000000000",
		266 =>	"00000001000000000000001000000010",
		267 =>	"00000010000000100000001000000010",
		268 =>	"00000001000000000000001000000010",
		269 =>	"00000010000000100000001000000010",
		270 =>	"00000001000000010000000100000001",
		271 =>	"00000001000000010000000100000001",
		272 =>	"00000011000000110000001100000011", -- IMG_8x8_BULLET
		273 =>	"00000011000000110000001100000011",
		274 =>	"00000011000000110000001100000011",
		275 =>	"00000011000000110000001100000011",
		276 =>	"00000011000000110000001100000100",
		277 =>	"00000011000000110000001100000011",
		278 =>	"00000011000000110000010000000100",
		279 =>	"00000100000000110000001100000011",
		280 =>	"00000011000000110000010000000100",
		281 =>	"00000100000000110000001100000011",
		282 =>	"00000011000000110000010000000100",
		283 =>	"00000100000000110000001100000011",
		284 =>	"00000011000000110000001100000011",
		285 =>	"00000011000000110000001100000011",
		286 =>	"00000011000000110000001100000011",
		287 =>	"00000011000000110000001100000011",
		288 =>	"00000011000001010000010100000101", -- IMG_8x8_GRASS
		289 =>	"00000110000001010000011100000011",
		290 =>	"00000101000001010000011000000111",
		291 =>	"00000101000001110000010100000111",
		292 =>	"00000101000001010000010100000101",
		293 =>	"00000101000001110000011100000111",
		294 =>	"00000110000001010000010100000111",
		295 =>	"00000111000001100000010100000111",
		296 =>	"00000101000001010000011100000110",
		297 =>	"00000111000001110000011100000110",
		298 =>	"00000101000001100000010100000111",
		299 =>	"00000111000001110000011100000111",
		300 =>	"00000111000001110000011100000111",
		301 =>	"00000111000001100000011100000111",
		302 =>	"00000011000001110000011100000110",
		303 =>	"00000111000001110000011100000011",
		304 =>	"00000001000001000000010000001000", -- IMG_8x8_ICE
		305 =>	"00000001000001000000010000001000",
		306 =>	"00000100000001000000010000000100",
		307 =>	"00000100000001000000100000000001",
		308 =>	"00000100000001000000010000000100",
		309 =>	"00000100000010000000000100000100",
		310 =>	"00001000000001000000010000000100",
		311 =>	"00001000000000010000010000000100",
		312 =>	"00000001000001000000010000001000",
		313 =>	"00000001000001000000010000001000",
		314 =>	"00000100000001000000100000000001",
		315 =>	"00000100000001000000100000000001",
		316 =>	"00000100000010000000000100000100",
		317 =>	"00000100000010000000000100000100",
		318 =>	"00001000000000010000010000000100",
		319 =>	"00001000000000010000010000000100",
		320 =>	"00000100000001000000010000000100", -- IMG_8x8_IRON
		321 =>	"00000100000001000000010000000100",
		322 =>	"00000100000001000000010000000100",
		323 =>	"00000100000001000000010000000001",
		324 =>	"00000100000001000000100000001000",
		325 =>	"00001000000010000000000100000001",
		326 =>	"00000100000001000000100000001000",
		327 =>	"00001000000010000000000100000001",
		328 =>	"00000100000001000000100000001000",
		329 =>	"00001000000010000000000100000001",
		330 =>	"00000100000001000000100000001000",
		331 =>	"00001000000010000000000100000001",
		332 =>	"00000100000001000000000100000001",
		333 =>	"00000001000000010000000100000001",
		334 =>	"00000100000000010000000100000001",
		335 =>	"00000001000000010000000100000001",
		336 =>	"00000001000000010000000100000010", -- IMG_8x8_LIVES_REMAINING_ICON
		337 =>	"00000010000000100000000100000001",
		338 =>	"00000001000000100000000100000001",
		339 =>	"00000010000000010000000100000010",
		340 =>	"00000001000000100000000100000010",
		341 =>	"00000010000000100000000100000010",
		342 =>	"00000001000000100000001000000010",
		343 =>	"00000001000000100000001000000010",
		344 =>	"00000001000000100000001000000001",
		345 =>	"00000001000000010000001000000010",
		346 =>	"00000001000000100000001000000010",
		347 =>	"00000001000000100000001000000010",
		348 =>	"00000001000000100000000100000010",
		349 =>	"00000010000000100000000100000010",
		350 =>	"00000001000000100000000100000001",
		351 =>	"00000010000000010000000100000010",
		352 =>	"00001001000010010000100100001001", -- IMG_8x8_NULL
		353 =>	"00001001000010010000100100001001",
		354 =>	"00001001000010010000100100001010",
		355 =>	"00001001000010010000100100001001",
		356 =>	"00001001000010010000101000001001",
		357 =>	"00001001000010010000100100001001",
		358 =>	"00001001000010010000100100001001",
		359 =>	"00001001000010010000100100001001",
		360 =>	"00001001000010010000101100001001",
		361 =>	"00001001000010010000100100001001",
		362 =>	"00001001000010010000100100001001",
		363 =>	"00001001000010010000100100001001",
		364 =>	"00001001000010010000100100001001",
		365 =>	"00001001000010010000100100001001",
		366 =>	"00001001000010010000100100001001",
		367 =>	"00001001000010010000100100001001",
		368 =>	"00000001000000010000000100000001", -- IMG_8x8_TANKS_REMAINING_ICON
		369 =>	"00000001000000010000000100000001",
		370 =>	"00000001000000110000000100000001",
		371 =>	"00000011000000010000000100000011",
		372 =>	"00000001000000110000000100000011",
		373 =>	"00000011000000110000000100000011",
		374 =>	"00000001000000110000001100000011",
		375 =>	"00000000000000110000001100000011",
		376 =>	"00000001000000110000001100000011",
		377 =>	"00000000000000110000001100000011",
		378 =>	"00000001000000110000000100000011",
		379 =>	"00000011000000110000000100000011",
		380 =>	"00000001000000110000000100000001",
		381 =>	"00000011000000010000000100000011",
		382 =>	"00000001000000010000000100000011",
		383 =>	"00000011000000110000000100000001",
		384 =>	"00001100000011000000110000001100", -- IMG_8x8_WATER
		385 =>	"00001100000011000000110000001101",
		386 =>	"00001100000011010000110000001100",
		387 =>	"00001100000011000000110000001100",
		388 =>	"00001100000011000000110100001100",
		389 =>	"00001100000011000000110000001100",
		390 =>	"00001100000011000000110000001101",
		391 =>	"00001100000011000000110100001100",
		392 =>	"00001100000011000000110000001100",
		393 =>	"00001100000011000000110000001101",
		394 =>	"00001100000011000000110000001101",
		395 =>	"00001100000011000000110000001100",
		396 =>	"00001100000011000000110100001100",
		397 =>	"00001101000011000000110000001100",
		398 =>	"00001101000011000000110000001100",
		399 =>	"00001100000011000000110000001100",


--			***** 16x16 IMAGES *****


		400 =>	"00000011000000110000001100000011", -- IMG_16x16_BASE_ALIVE
		401 =>	"00000011000000110000001100000011",
		402 =>	"00000011000000110000001100000011",
		403 =>	"00000011000000110000001100000011",
		404 =>	"00000001000000010000001100000011",
		405 =>	"00000011000000110000001100000011",
		406 =>	"00000011000000110000001100000011",
		407 =>	"00000011000000110000000100000001",
		408 =>	"00000011000000010000000100000011",
		409 =>	"00000011000000110000000100000001",
		410 =>	"00000001000000110000001100000011",
		411 =>	"00000011000000010000000100000011",
		412 =>	"00000001000000010000000100000001",
		413 =>	"00000011000000110000001100000001",
		414 =>	"00000000000000010000001100000011",
		415 =>	"00000001000000010000000100000001",
		416 =>	"00000011000000010000000100000001",
		417 =>	"00000011000000110000001100000001",
		418 =>	"00000001000000110000001100000011",
		419 =>	"00000001000000010000000100000011",
		420 =>	"00000001000000010000000100000001",
		421 =>	"00000001000000010000001100000001",
		422 =>	"00000001000000110000000100000001",
		423 =>	"00000001000000010000000100000001",
		424 =>	"00000011000000110000000100000000",
		425 =>	"00000001000000010000000100000001",
		426 =>	"00000001000000010000000100000001",
		427 =>	"00000000000000010000001100000011",
		428 =>	"00000011000000010000000100000001",
		429 =>	"00000000000000010000000100000001",
		430 =>	"00000001000000010000000100000000",
		431 =>	"00000001000000010000000100000011",
		432 =>	"00000011000000110000000100000001",
		433 =>	"00000001000000010000000000000001",
		434 =>	"00000001000000000000000100000001",
		435 =>	"00000001000000010000001100000011",
		436 =>	"00000011000000110000000100000001",
		437 =>	"00000001000000010000000100000001",
		438 =>	"00000001000000010000000100000001",
		439 =>	"00000001000000010000001100000011",
		440 =>	"00000011000000110000001100000001",
		441 =>	"00000001000000010000001100000001",
		442 =>	"00000001000000110000000100000001",
		443 =>	"00000001000000110000001100000011",
		444 =>	"00000011000000110000001100000011",
		445 =>	"00000011000000110000001100000001",
		446 =>	"00000001000000110000001100000011",
		447 =>	"00000011000000110000001100000011",
		448 =>	"00000011000000110000001100000011",
		449 =>	"00000011000000110000000100000001",
		450 =>	"00000001000000010000001100000011",
		451 =>	"00000011000000110000001100000011",
		452 =>	"00000011000000110000001100000011",
		453 =>	"00000001000000010000000100000001",
		454 =>	"00000001000000010000000100000001",
		455 =>	"00000011000000110000001100000011",
		456 =>	"00000011000000110000001100000011",
		457 =>	"00000001000000010000001100000001",
		458 =>	"00000001000000110000000100000001",
		459 =>	"00000011000000110000001100000011",
		460 =>	"00000011000000110000001100000011",
		461 =>	"00000011000000110000001100000011",
		462 =>	"00000011000000110000001100000011",
		463 =>	"00000011000000110000001100000011",
		464 =>	"00000011000000110000001100000011", -- IMG_16x16_BASE_DEAD
		465 =>	"00000011000000110000001100000011",
		466 =>	"00000011000000110000001100000011",
		467 =>	"00000011000000110000001100000011",
		468 =>	"00000011000000110000001100000011",
		469 =>	"00000011000000100000001100000011",
		470 =>	"00000011000000110000001100000011",
		471 =>	"00000011000000110000001100000011",
		472 =>	"00000011000000110000001100000011",
		473 =>	"00000010000000100000001100000001",
		474 =>	"00000011000000110000001100000011",
		475 =>	"00000011000000110000001100000011",
		476 =>	"00000011000000110000001100000011",
		477 =>	"00000010000000110000000100000001",
		478 =>	"00000001000000110000001100000011",
		479 =>	"00000011000000110000001100000011",
		480 =>	"00000011000000110000001100000010",
		481 =>	"00000011000000010000000100000001",
		482 =>	"00000001000000010000001100000011",
		483 =>	"00000011000000110000001100000011",
		484 =>	"00000011000000110000001000000010",
		485 =>	"00000011000000010000000100000001",
		486 =>	"00000001000000010000000100000001",
		487 =>	"00000001000000110000001100000011",
		488 =>	"00000011000000110000001000000011",
		489 =>	"00000001000000010000000100000001",
		490 =>	"00000001000000010000000100000001",
		491 =>	"00000001000000010000001100000011",
		492 =>	"00000011000000100000001000000011",
		493 =>	"00000001000000010000000100000001",
		494 =>	"00000001000000010000000100000001",
		495 =>	"00000001000000010000001100000011",
		496 =>	"00000011000000100000001100000011",
		497 =>	"00000001000000010000000100000001",
		498 =>	"00000001000000010000000100000001",
		499 =>	"00000011000000010000000100000011",
		500 =>	"00000011000000100000001100000001",
		501 =>	"00000001000000010000000100000001",
		502 =>	"00000001000000110000001100000001",
		503 =>	"00000011000000010000000100000011",
		504 =>	"00000011000000100000001100000011",
		505 =>	"00000011000000010000000100000001",
		506 =>	"00000011000000110000001100000011",
		507 =>	"00000011000000010000001100000011",
		508 =>	"00000011000000100000001100000011",
		509 =>	"00000011000000110000001100000001",
		510 =>	"00000011000000110000001100000011",
		511 =>	"00000011000000010000001100000011",
		512 =>	"00000011000000100000001100000011",
		513 =>	"00000011000000110000001100000011",
		514 =>	"00000011000000110000001100000011",
		515 =>	"00000011000000110000001100000011",
		516 =>	"00000011000000100000001100000011",
		517 =>	"00000011000000110000001100000011",
		518 =>	"00000011000000110000001100000011",
		519 =>	"00000011000000110000001100000011",
		520 =>	"00000011000000100000001100000011",
		521 =>	"00000011000000110000001100000011",
		522 =>	"00000011000000110000001100000011",
		523 =>	"00000011000000110000001100000011",
		524 =>	"00000011000000110000001100000011",
		525 =>	"00000011000000110000001100000011",
		526 =>	"00000011000000110000001100000011",
		527 =>	"00000011000000110000001100000011",
		528 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_BOMB
		529 =>	"00000011000000110000001100000011",
		530 =>	"00000011000000110000001100000011",
		531 =>	"00000011000000110000001100000011",
		532 =>	"00000011000010000000100000001000",
		533 =>	"00001000000010000000100000001000",
		534 =>	"00001000000010000000100000001000",
		535 =>	"00001000000010000000010000000011",
		536 =>	"00001000000000110000001100000011",
		537 =>	"00000011000000110000001100000011",
		538 =>	"00000011000000110000001100000011",
		539 =>	"00000011000000110000100000001110",
		540 =>	"00001000000000110000111000001110",
		541 =>	"00001110000010000000100000001000",
		542 =>	"00000100000001000000001100001110",
		543 =>	"00001110000011100000100000001110",
		544 =>	"00001000000000110000111000001110",
		545 =>	"00001110000010000000010000001110",
		546 =>	"00000011000000110000010000000011",
		547 =>	"00001110000011100000100000001110",
		548 =>	"00001000000000110000111000001110",
		549 =>	"00001000000001000000010000000100",
		550 =>	"00001110000000110000001100000100",
		551 =>	"00000011000011100000100000001110",
		552 =>	"00001000000000110000111000001000",
		553 =>	"00000100000011100000100000000100",
		554 =>	"00001110000001000000001100000100",
		555 =>	"00000011000011100000100000001110",
		556 =>	"00001000000000110000111000000100",
		557 =>	"00000011000001000000001100000011",
		558 =>	"00000100000000110000001100000100",
		559 =>	"00000011000011100000100000001110",
		560 =>	"00001000000000110000111000001000",
		561 =>	"00000100000011100000100000000100",
		562 =>	"00001110000001000000001100000100",
		563 =>	"00000011000011100000100000001110",
		564 =>	"00001000000000110000111000000100",
		565 =>	"00000011000001000000001100000011",
		566 =>	"00000100000000110000001100000100",
		567 =>	"00000011000011100000100000001110",
		568 =>	"00001000000000110000111000001000",
		569 =>	"00000100000011100000100000000100",
		570 =>	"00001110000001000000001100000011",
		571 =>	"00001110000011100000100000001110",
		572 =>	"00001000000000110000111000001110",
		573 =>	"00000100000011100000001100000011",
		574 =>	"00000100000000110000111000001110",
		575 =>	"00001110000011100000100000001110",
		576 =>	"00001000000000110000111000001110",
		577 =>	"00001110000010000000010000000100",
		578 =>	"00000011000011100000111000001110",
		579 =>	"00001110000011100000100000001110",
		580 =>	"00001000000000110000111000001110",
		581 =>	"00001110000000110000001100000011",
		582 =>	"00001110000011100000111000001110",
		583 =>	"00001110000011100000100000001110",
		584 =>	"00000100000010000000100000001000",
		585 =>	"00001000000010000000100000001000",
		586 =>	"00001000000010000000100000001000",
		587 =>	"00001000000010000000010000001110",
		588 =>	"00000011000011100000111000001110",
		589 =>	"00001110000011100000111000001110",
		590 =>	"00001110000011100000111000001110",
		591 =>	"00001110000011100000111000000011",
		592 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_GUN
		593 =>	"00000011000000110000001100000011",
		594 =>	"00000011000000110000001100000011",
		595 =>	"00000011000000110000001100000011",
		596 =>	"00000011000010000000100000001000",
		597 =>	"00001000000010000000100000001000",
		598 =>	"00001000000010000000100000001000",
		599 =>	"00001000000010000000010000000011",
		600 =>	"00001000000000110000001100000011",
		601 =>	"00000011000000110000001100000011",
		602 =>	"00000011000000110000001100000011",
		603 =>	"00000011000000110000100000001110",
		604 =>	"00001000000000110000111000001110",
		605 =>	"00001110000011100000111000001110",
		606 =>	"00001110000011100000111000001110",
		607 =>	"00001110000011100000100000001110",
		608 =>	"00001000000000110000111000001000",
		609 =>	"00001110000011100000111000001110",
		610 =>	"00001110000011100000111000001110",
		611 =>	"00001110000011100000100000001110",
		612 =>	"00001000000000110000010000001000",
		613 =>	"00001000000010000000100000001000",
		614 =>	"00001000000010000000010000000011",
		615 =>	"00001110000011100000100000001110",
		616 =>	"00001000000000110000100000000100",
		617 =>	"00000100000001000000010000000100",
		618 =>	"00000100000001000000010000000100",
		619 =>	"00000011000011100000100000001110",
		620 =>	"00001000000000110000001100000100",
		621 =>	"00000100000011100000111000001110",
		622 =>	"00001110000011100000111000000100",
		623 =>	"00000011000011100000100000001110",
		624 =>	"00001000000000110000111000000011",
		625 =>	"00000011000001000000010000001110",
		626 =>	"00000100000001000000010000000100",
		627 =>	"00000100000000110000100000001110",
		628 =>	"00001000000000110000111000001110",
		629 =>	"00001110000000110000010000000011",
		630 =>	"00000011000001000000100000001110",
		631 =>	"00000100000000110000100000001110",
		632 =>	"00001000000000110000111000001110",
		633 =>	"00001110000011100000001100000100",
		634 =>	"00000100000001000000100000001110",
		635 =>	"00000100000000110000100000001110",
		636 =>	"00001000000000110000111000001110",
		637 =>	"00001110000011100000111000000011",
		638 =>	"00000011000001000000111000001110",
		639 =>	"00000100000000110000100000001110",
		640 =>	"00001000000000110000111000001110",
		641 =>	"00001110000011100000111000001110",
		642 =>	"00001110000001000000010000000100",
		643 =>	"00000100000000110000100000001110",
		644 =>	"00001000000000110000111000001110",
		645 =>	"00001110000011100000111000001110",
		646 =>	"00001110000000110000001100000011",
		647 =>	"00000011000011100000100000001110",
		648 =>	"00000100000010000000100000001000",
		649 =>	"00001000000010000000100000001000",
		650 =>	"00001000000010000000100000001000",
		651 =>	"00001000000010000000010000001110",
		652 =>	"00000011000011100000111000001110",
		653 =>	"00001110000011100000111000001110",
		654 =>	"00001110000011100000111000001110",
		655 =>	"00001110000011100000111000000011",
		656 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_SHELL
		657 =>	"00000011000000110000001100000011",
		658 =>	"00000011000000110000001100000011",
		659 =>	"00000011000000110000001100000011",
		660 =>	"00000011000010000000100000001000",
		661 =>	"00001000000010000000100000001000",
		662 =>	"00001000000010000000100000001000",
		663 =>	"00001000000010000000010000000011",
		664 =>	"00001000000000110000001100000011",
		665 =>	"00000011000000110000001100000011",
		666 =>	"00000011000000110000001100000011",
		667 =>	"00000011000000110000100000001110",
		668 =>	"00001000000000110000111000001110",
		669 =>	"00001110000011100000111000001110",
		670 =>	"00001110000011100000111000001110",
		671 =>	"00001110000011100000100000001110",
		672 =>	"00001000000000110000111000001110",
		673 =>	"00001110000011100000111000001110",
		674 =>	"00001110000011100000111000001110",
		675 =>	"00001110000011100000100000001110",
		676 =>	"00001000000000110000111000001110",
		677 =>	"00001110000010000000100000001000",
		678 =>	"00000100000001000000001100001110",
		679 =>	"00001110000011100000100000001110",
		680 =>	"00001000000000110000111000001110",
		681 =>	"00001000000010000000010000000100",
		682 =>	"00000100000001000000010000000011",
		683 =>	"00001110000011100000100000001110",
		684 =>	"00001000000000110000111000001110",
		685 =>	"00001000000001000000010000000100",
		686 =>	"00000100000001000000010000000011",
		687 =>	"00001110000011100000100000001110",
		688 =>	"00001000000000110000111000001110",
		689 =>	"00000100000001000000010000000100",
		690 =>	"00000100000001000000010000000011",
		691 =>	"00001110000011100000100000001110",
		692 =>	"00001000000000110000111000000100",
		693 =>	"00000100000001000000010000000100",
		694 =>	"00000100000001000000010000000011",
		695 =>	"00001110000011100000100000001110",
		696 =>	"00001000000000110000111000000011",
		697 =>	"00000011000000110000001100000011",
		698 =>	"00000100000001000000010000000100",
		699 =>	"00000011000011100000100000001110",
		700 =>	"00001000000000110000111000001110",
		701 =>	"00001110000011100000111000001110",
		702 =>	"00000011000000110000001100000011",
		703 =>	"00000011000011100000100000001110",
		704 =>	"00001000000000110000111000001110",
		705 =>	"00001110000011100000111000001110",
		706 =>	"00001110000011100000111000001110",
		707 =>	"00001110000011100000100000001110",
		708 =>	"00001000000000110000111000001110",
		709 =>	"00001110000011100000111000001110",
		710 =>	"00001110000011100000111000001110",
		711 =>	"00001110000011100000100000001110",
		712 =>	"00000100000010000000100000001000",
		713 =>	"00001000000010000000100000001000",
		714 =>	"00001000000010000000100000001000",
		715 =>	"00001000000010000000010000001110",
		716 =>	"00000011000011100000111000001110",
		717 =>	"00001110000011100000111000001110",
		718 =>	"00001110000011100000111000001110",
		719 =>	"00001110000011100000111000000011",
		720 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_SHOVEL
		721 =>	"00000011000000110000001100000011",
		722 =>	"00000011000000110000001100000011",
		723 =>	"00000011000000110000001100000011",
		724 =>	"00000011000010000000100000001000",
		725 =>	"00001000000010000000100000001000",
		726 =>	"00001000000010000000100000001000",
		727 =>	"00001000000010000000010000000011",
		728 =>	"00001000000000110000001100000011",
		729 =>	"00000011000000110000001100000011",
		730 =>	"00000011000000110000001100000011",
		731 =>	"00000011000000110000100000001110",
		732 =>	"00001000000000110000111000001110",
		733 =>	"00001110000011100000111000001110",
		734 =>	"00001110000011100000100000001110",
		735 =>	"00001110000011100000100000001110",
		736 =>	"00001000000000110000111000001110",
		737 =>	"00001110000011100000111000001110",
		738 =>	"00001110000011100000100000000100",
		739 =>	"00001110000011100000100000001110",
		740 =>	"00001000000000110000111000001110",
		741 =>	"00001110000011100000111000001110",
		742 =>	"00001110000011100000010000000100",
		743 =>	"00000100000011100000100000001110",
		744 =>	"00001000000000110000111000001110",
		745 =>	"00001110000011100000111000001110",
		746 =>	"00001110000010000000001100000011",
		747 =>	"00000011000011100000100000001110",
		748 =>	"00001000000000110000111000001110",
		749 =>	"00001110000010000000111000001110",
		750 =>	"00001000000000110000111000001110",
		751 =>	"00001110000011100000100000001110",
		752 =>	"00001000000000110000111000001110",
		753 =>	"00001000000010000000010000001000",
		754 =>	"00000011000011100000111000001110",
		755 =>	"00001110000011100000100000001110",
		756 =>	"00001000000000110000111000001000",
		757 =>	"00001000000001000000111000000100",
		758 =>	"00000011000011100000111000001110",
		759 =>	"00001110000011100000100000001110",
		760 =>	"00001000000000110000111000001000",
		761 =>	"00000100000011100000010000000100",
		762 =>	"00000100000000110000111000001110",
		763 =>	"00001110000011100000100000001110",
		764 =>	"00001000000000110000111000000100",
		765 =>	"00000100000001000000010000000100",
		766 =>	"00000011000011100000111000001110",
		767 =>	"00001110000011100000100000001110",
		768 =>	"00001000000000110000111000000100",
		769 =>	"00000100000001000000010000000011",
		770 =>	"00001110000011100000111000001110",
		771 =>	"00001110000011100000100000001110",
		772 =>	"00001000000000110000111000000011",
		773 =>	"00000011000000110000001100001110",
		774 =>	"00001110000011100000111000001110",
		775 =>	"00001110000011100000100000001110",
		776 =>	"00000100000010000000100000001000",
		777 =>	"00001000000010000000100000001000",
		778 =>	"00001000000010000000100000001000",
		779 =>	"00001000000010000000010000001110",
		780 =>	"00000011000011100000111000001110",
		781 =>	"00001110000011100000111000001110",
		782 =>	"00001110000011100000111000001110",
		783 =>	"00001110000011100000111000000011",
		784 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_STAR
		785 =>	"00000011000000110000001100000011",
		786 =>	"00000011000000110000001100000011",
		787 =>	"00000011000000110000001100000011",
		788 =>	"00000011000010000000100000001000",
		789 =>	"00001000000010000000100000001000",
		790 =>	"00001000000010000000100000001000",
		791 =>	"00001000000010000000010000000011",
		792 =>	"00001000000000110000001100000011",
		793 =>	"00000011000000110000001100000011",
		794 =>	"00000011000000110000001100000011",
		795 =>	"00000011000000110000100000001110",
		796 =>	"00001000000000110000111000001110",
		797 =>	"00001110000011100000111000001000",
		798 =>	"00000011000011100000111000001110",
		799 =>	"00001110000011100000100000001110",
		800 =>	"00001000000000110000111000001110",
		801 =>	"00001110000011100000100000001000",
		802 =>	"00000100000000110000111000001110",
		803 =>	"00001110000011100000100000001110",
		804 =>	"00001000000000110000111000001110",
		805 =>	"00001110000011100000100000001000",
		806 =>	"00000100000000110000111000001110",
		807 =>	"00001110000011100000100000001110",
		808 =>	"00001000000000110000100000001000",
		809 =>	"00001000000010000000100000000100",
		810 =>	"00000100000010000000100000001000",
		811 =>	"00001000000000110000100000001110",
		812 =>	"00001000000000110000111000000100",
		813 =>	"00000100000001000000100000000100",
		814 =>	"00001000000001000000010000000100",
		815 =>	"00000011000000110000100000001110",
		816 =>	"00001000000000110000111000001110",
		817 =>	"00000100000010000000100000001000",
		818 =>	"00001000000001000000010000000011",
		819 =>	"00000011000011100000100000001110",
		820 =>	"00001000000000110000111000001110",
		821 =>	"00001000000010000000010000000100",
		822 =>	"00001000000010000000010000000011",
		823 =>	"00001110000011100000100000001110",
		824 =>	"00001000000000110000111000000100",
		825 =>	"00001000000001000000010000000011",
		826 =>	"00000100000001000000100000000100",
		827 =>	"00000011000011100000100000001110",
		828 =>	"00001000000000110000111000001000",
		829 =>	"00000100000001000000001100000011",
		830 =>	"00000011000001000000010000001000",
		831 =>	"00000011000011100000100000001110",
		832 =>	"00001000000000110000111000000100",
		833 =>	"00000011000000110000001100001110",
		834 =>	"00001110000000110000001100000100",
		835 =>	"00000011000011100000100000001110",
		836 =>	"00001000000000110000111000000011",
		837 =>	"00000011000011100000111000001110",
		838 =>	"00001110000011100000111000000011",
		839 =>	"00000011000011100000100000001110",
		840 =>	"00000100000010000000100000001000",
		841 =>	"00001000000010000000100000001000",
		842 =>	"00001000000010000000100000001000",
		843 =>	"00001000000010000000010000001110",
		844 =>	"00000011000011100000111000001110",
		845 =>	"00001110000011100000111000001110",
		846 =>	"00001110000011100000111000001110",
		847 =>	"00001110000011100000111000000011",
		848 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_TANK
		849 =>	"00000011000000110000001100000011",
		850 =>	"00000011000000110000001100000011",
		851 =>	"00000011000000110000001100000011",
		852 =>	"00000011000010000000100000001000",
		853 =>	"00001000000010000000100000001000",
		854 =>	"00001000000010000000100000001000",
		855 =>	"00001000000010000000010000000011",
		856 =>	"00001000000000110000001100000011",
		857 =>	"00000011000000110000001100000011",
		858 =>	"00000011000000110000001100000011",
		859 =>	"00000011000000110000100000001110",
		860 =>	"00001000000000110000111000001110",
		861 =>	"00001110000011100000111000001110",
		862 =>	"00001110000011100000111000001110",
		863 =>	"00001110000011100000100000001110",
		864 =>	"00001000000000110000111000001000",
		865 =>	"00001110000011100000111000001110",
		866 =>	"00001110000011100000111000001110",
		867 =>	"00001110000011100000100000001110",
		868 =>	"00001000000000110000010000001000",
		869 =>	"00001000000010000000100000001000",
		870 =>	"00001000000010000000010000000011",
		871 =>	"00001110000011100000100000001110",
		872 =>	"00001000000000110000100000000100",
		873 =>	"00000100000001000000010000000100",
		874 =>	"00000100000001000000010000000100",
		875 =>	"00000011000011100000100000001110",
		876 =>	"00001000000000110000001100000100",
		877 =>	"00000100000011100000111000001110",
		878 =>	"00001110000011100000111000000100",
		879 =>	"00000011000011100000100000001110",
		880 =>	"00001000000000110000111000000011",
		881 =>	"00000011000001000000010000001110",
		882 =>	"00000100000001000000010000000100",
		883 =>	"00000100000000110000100000001110",
		884 =>	"00001000000000110000111000001110",
		885 =>	"00001110000000110000010000000011",
		886 =>	"00000011000001000000100000001110",
		887 =>	"00000100000000110000100000001110",
		888 =>	"00001000000000110000111000001110",
		889 =>	"00001110000011100000001100000100",
		890 =>	"00000100000001000000100000001110",
		891 =>	"00000100000000110000100000001110",
		892 =>	"00001000000000110000111000001110",
		893 =>	"00001110000011100000111000000011",
		894 =>	"00000011000001000000111000001110",
		895 =>	"00000100000000110000100000001110",
		896 =>	"00001000000000110000111000001110",
		897 =>	"00001110000011100000111000001110",
		898 =>	"00001110000001000000010000000100",
		899 =>	"00000100000000110000100000001110",
		900 =>	"00001000000000110000111000001110",
		901 =>	"00001110000011100000111000001110",
		902 =>	"00001110000000110000001100000011",
		903 =>	"00000011000011100000100000001110",
		904 =>	"00000100000010000000100000001000",
		905 =>	"00001000000010000000100000001000",
		906 =>	"00001000000010000000100000001000",
		907 =>	"00001000000010000000010000001110",
		908 =>	"00000011000011100000111000001110",
		909 =>	"00001110000011100000111000001110",
		910 =>	"00001110000011100000111000001110",
		911 =>	"00001110000011100000111000000011",
		912 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_TIME
		913 =>	"00000011000000110000001100000011",
		914 =>	"00000011000000110000001100000011",
		915 =>	"00000011000000110000001100000011",
		916 =>	"00000011000000110000100000001000",
		917 =>	"00001000000010000000100000001000",
		918 =>	"00001000000010000000100000001000",
		919 =>	"00001000000010000000100000000100",
		920 =>	"00001110000010000000001100000011",
		921 =>	"00000011000000110000001100000011",
		922 =>	"00000011000000110000001100000011",
		923 =>	"00000011000000110000001100001000",
		924 =>	"00001110000010000000001100001110",
		925 =>	"00001110000011100000111000001000",
		926 =>	"00000100000010000000010000000011",
		927 =>	"00001110000011100000111000001000",
		928 =>	"00001110000010000000001100001110",
		929 =>	"00001110000011100000111000000100",
		930 =>	"00000011000000110000001100001000",
		931 =>	"00000100000000110000111000001000",
		932 =>	"00001110000010000000001100001110",
		933 =>	"00001110000011100000010000000100",
		934 =>	"00000100000001000000001100000011",
		935 =>	"00000011000000110000111000001000",
		936 =>	"00001110000010000000001100001110",
		937 =>	"00001110000001000000100000001000",
		938 =>	"00001000000010000000010000000011",
		939 =>	"00001110000011100000111000001000",
		940 =>	"00001110000010000000001100001110",
		941 =>	"00000100000010000000100000001110",
		942 =>	"00001000000010000000100000000100",
		943 =>	"00000011000011100000111000001000",
		944 =>	"00001110000010000000001100001110",
		945 =>	"00000100000010000000100000001110",
		946 =>	"00001000000010000000100000000100",
		947 =>	"00000011000011100000111000001000",
		948 =>	"00001110000010000000001100001110",
		949 =>	"00000100000010000000100000001000",
		950 =>	"00001110000010000000100000000100",
		951 =>	"00000011000011100000111000001000",
		952 =>	"00001110000010000000001100001110",
		953 =>	"00000011000001000000100000001000",
		954 =>	"00001000000010000000010000000011",
		955 =>	"00001110000011100000111000001000",
		956 =>	"00001110000010000000001100001110",
		957 =>	"00001110000000110000010000000100",
		958 =>	"00000100000001000000001100001110",
		959 =>	"00001110000011100000111000001000",
		960 =>	"00001110000010000000001100001110",
		961 =>	"00001110000011100000001100000011",
		962 =>	"00000011000000110000111000001110",
		963 =>	"00001110000011100000111000001000",
		964 =>	"00001110000010000000001100001110",
		965 =>	"00001110000011100000111000001110",
		966 =>	"00001110000011100000111000001110",
		967 =>	"00001110000011100000111000001000",
		968 =>	"00001110000001000000100000001000",
		969 =>	"00001000000010000000100000001000",
		970 =>	"00001000000010000000100000001000",
		971 =>	"00001000000010000000100000000100",
		972 =>	"00000011000000110000111000001110",
		973 =>	"00001110000011100000111000001110",
		974 =>	"00001110000011100000111000001110",
		975 =>	"00001110000011100000111000001110",
		976 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK1
		977 =>	"00000011000000110000001100000011",
		978 =>	"00000011000000110000001100000011",
		979 =>	"00000011000000110000001100000011",
		980 =>	"00000011000000110000001100000011",
		981 =>	"00000011000000110000001100001000",
		982 =>	"00000011000000110000001100000011",
		983 =>	"00000011000000110000001100000011",
		984 =>	"00000011000000110000001100000011",
		985 =>	"00000011000000110000001100001000",
		986 =>	"00000011000000110000001100000011",
		987 =>	"00000011000000110000001100000011",
		988 =>	"00000011000000110000001100000011",
		989 =>	"00000011000000110000001100001000",
		990 =>	"00000011000000110000001100000011",
		991 =>	"00000011000000110000001100000011",
		992 =>	"00000011000010000000010000000100",
		993 =>	"00000011000000110000010000001000",
		994 =>	"00001110000000110000001100001000",
		995 =>	"00000100000001000000001100000011",
		996 =>	"00000011000011100000111000000100",
		997 =>	"00000011000010000000010000001000",
		998 =>	"00001110000011100000001100000100",
		999 =>	"00001110000011100000001100000011",
		1000 =>	"00000011000010000000010000000100",
		1001 =>	"00001000000010000000010000001000",
		1002 =>	"00001110000011100000111000000100",
		1003 =>	"00000100000001000000001100000011",
		1004 =>	"00000011000011100000111000000100",
		1005 =>	"00001000000010000000010000000100",
		1006 =>	"00000100000011100000111000000100",
		1007 =>	"00001110000011100000001100000011",
		1008 =>	"00000011000010000000010000000100",
		1009 =>	"00001000000001000000010000001110",
		1010 =>	"00000100000001000000111000000100",
		1011 =>	"00000100000001000000001100000011",
		1012 =>	"00000011000011100000111000000100",
		1013 =>	"00001000000001000000111000001110",
		1014 =>	"00001000000001000000111000000100",
		1015 =>	"00001110000011100000001100000011",
		1016 =>	"00000011000010000000010000000100",
		1017 =>	"00001000000001000000111000001000",
		1018 =>	"00001000000001000000111000000100",
		1019 =>	"00000100000001000000001100000011",
		1020 =>	"00000011000011100000111000000100",
		1021 =>	"00001000000001000000010000000100",
		1022 =>	"00000100000001000000111000000100",
		1023 =>	"00001110000011100000001100000011",
		1024 =>	"00000011000010000000010000000100",
		1025 =>	"00001000000010000000010000000100",
		1026 =>	"00000100000011100000111000000100",
		1027 =>	"00000100000001000000001100000011",
		1028 =>	"00000011000011100000111000000100",
		1029 =>	"00000011000010000000010000000100",
		1030 =>	"00001110000011100000001100000100",
		1031 =>	"00001110000011100000001100000011",
		1032 =>	"00000011000010000000010000000100",
		1033 =>	"00000011000000110000111000001110",
		1034 =>	"00001110000000110000001100000100",
		1035 =>	"00000100000001000000001100000011",
		1036 =>	"00000011000000110000001100000011",
		1037 =>	"00000011000000110000001100000100",
		1038 =>	"00000011000000110000001100000011",
		1039 =>	"00000011000000110000001100000011",
		1040 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK2
		1041 =>	"00000011000000110000001100000011",
		1042 =>	"00000011000000110000001100000011",
		1043 =>	"00000011000000110000001100000011",
		1044 =>	"00000011000000110000001100000011",
		1045 =>	"00000011000000110000001100001000",
		1046 =>	"00000011000000110000001100000011",
		1047 =>	"00000011000000110000001100000011",
		1048 =>	"00000011000000110000001100000011",
		1049 =>	"00000011000000110000001100001000",
		1050 =>	"00000011000000110000001100000011",
		1051 =>	"00000011000000110000001100000011",
		1052 =>	"00000011000001000000111000000011",
		1053 =>	"00001000000010000000111000001000",
		1054 =>	"00001110000001000000010000000011",
		1055 =>	"00000100000011100000001100000011",
		1056 =>	"00000011000011100000111000001000",
		1057 =>	"00001000000010000000111000001000",
		1058 =>	"00001110000001000000010000000100",
		1059 =>	"00001110000011100000001100000011",
		1060 =>	"00000011000011100000111000000100",
		1061 =>	"00001000000010000000111000001000",
		1062 =>	"00001110000011100000111000000100",
		1063 =>	"00001110000011100000001100000011",
		1064 =>	"00000011000000110000001100000100",
		1065 =>	"00000100000010000000010000001000",
		1066 =>	"00000100000011100000111000000100",
		1067 =>	"00000011000000110000001100000011",
		1068 =>	"00000011000000110000001100000100",
		1069 =>	"00001000000001000000010000000100",
		1070 =>	"00000100000001000000111000000100",
		1071 =>	"00000011000000110000001100000011",
		1072 =>	"00000011000001000000111000000100",
		1073 =>	"00001000000001000000010000001110",
		1074 =>	"00000100000001000000111000000100",
		1075 =>	"00000100000011100000001100000011",
		1076 =>	"00000011000011100000111000000100",
		1077 =>	"00001000000001000000111000001110",
		1078 =>	"00001000000001000000111000000100",
		1079 =>	"00001110000011100000001100000011",
		1080 =>	"00000011000011100000111000000100",
		1081 =>	"00001000000001000000111000001000",
		1082 =>	"00001000000001000000111000000100",
		1083 =>	"00001110000011100000001100000011",
		1084 =>	"00000011000000110000001100000100",
		1085 =>	"00001000000001000000010000000100",
		1086 =>	"00000100000001000000111000000100",
		1087 =>	"00000011000000110000001100000011",
		1088 =>	"00000011000000110000001100000100",
		1089 =>	"00001000000010000000010000000100",
		1090 =>	"00000100000010000000111000000100",
		1091 =>	"00000011000000110000001100000011",
		1092 =>	"00000011000001000000111000000100",
		1093 =>	"00000100000001000000100000001000",
		1094 =>	"00001000000011100000111000000100",
		1095 =>	"00000100000011100000001100000011",
		1096 =>	"00000011000011100000111000000100",
		1097 =>	"00001110000011100000111000001110",
		1098 =>	"00001110000011100000111000000100",
		1099 =>	"00001110000011100000001100000011",
		1100 =>	"00000011000011100000111000000011",
		1101 =>	"00001110000011100000111000001000",
		1102 =>	"00001110000011100000111000000011",
		1103 =>	"00001110000011100000001100000011",
		1104 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK3
		1105 =>	"00000011000000110000001100000011",
		1106 =>	"00000011000000110000001100000011",
		1107 =>	"00000011000000110000001100000011",
		1108 =>	"00000011000000110000001100000011",
		1109 =>	"00000011000000110000100000001000",
		1110 =>	"00000100000000110000001100000011",
		1111 =>	"00000011000000110000001100000011",
		1112 =>	"00000011000000110000001100000011",
		1113 =>	"00000011000000110000001100001000",
		1114 =>	"00000011000000110000001100000011",
		1115 =>	"00000011000000110000001100000011",
		1116 =>	"00000011000000110000001100000011",
		1117 =>	"00000011000000110000001100001000",
		1118 =>	"00000011000000110000001100000011",
		1119 =>	"00000011000000110000001100000011",
		1120 =>	"00000011000010000000010000000100",
		1121 =>	"00000011000000110000010000001000",
		1122 =>	"00001110000000110000001100001000",
		1123 =>	"00000100000001000000001100000011",
		1124 =>	"00000011000011100000111000000100",
		1125 =>	"00000011000010000000010000001000",
		1126 =>	"00001110000011100000001100000100",
		1127 =>	"00001110000011100000001100000011",
		1128 =>	"00000011000010000000010000000100",
		1129 =>	"00001000000010000000010000001000",
		1130 =>	"00001110000011100000111000000100",
		1131 =>	"00000100000001000000001100000011",
		1132 =>	"00000011000011100000111000000100",
		1133 =>	"00001000000010000000010000000100",
		1134 =>	"00000100000011100000111000000100",
		1135 =>	"00001110000011100000001100000011",
		1136 =>	"00000011000010000000010000000100",
		1137 =>	"00001000000001000000010000001110",
		1138 =>	"00000100000001000000111000000100",
		1139 =>	"00000100000001000000001100000011",
		1140 =>	"00000011000011100000111000000100",
		1141 =>	"00001000000001000000111000001110",
		1142 =>	"00001000000001000000111000000100",
		1143 =>	"00001110000011100000001100000011",
		1144 =>	"00000011000010000000010000000100",
		1145 =>	"00001000000001000000111000001000",
		1146 =>	"00001000000001000000111000000100",
		1147 =>	"00000100000001000000001100000011",
		1148 =>	"00000011000011100000111000000100",
		1149 =>	"00001000000001000000010000000100",
		1150 =>	"00000100000001000000111000000100",
		1151 =>	"00001110000011100000001100000011",
		1152 =>	"00000011000010000000010000000100",
		1153 =>	"00001000000010000000010000000100",
		1154 =>	"00000100000011100000111000000100",
		1155 =>	"00000100000001000000001100000011",
		1156 =>	"00000011000011100000111000000100",
		1157 =>	"00000011000010000000100000000100",
		1158 =>	"00001110000011100000001100000100",
		1159 =>	"00001110000011100000001100000011",
		1160 =>	"00000011000010000000010000000100",
		1161 =>	"00000011000010000000100000001110",
		1162 =>	"00001110000011100000001100000100",
		1163 =>	"00000100000001000000001100000011",
		1164 =>	"00000011000011100000111000000100",
		1165 =>	"00000011000000110000010000001000",
		1166 =>	"00001110000000110000001100000100",
		1167 =>	"00001110000011100000001100000011",
		1168 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK4
		1169 =>	"00000011000000110000001100000011",
		1170 =>	"00000011000000110000001100000011",
		1171 =>	"00000011000000110000001100000011",
		1172 =>	"00000011000010000000010000000100",
		1173 =>	"00000011000000110000100000001000",
		1174 =>	"00000100000000110000001100001000",
		1175 =>	"00000100000001000000001100000011",
		1176 =>	"00000011000011100000111000000100",
		1177 =>	"00000100000011100000100000001000",
		1178 =>	"00000100000011100000010000000100",
		1179 =>	"00001110000011100000001100000011",
		1180 =>	"00000011000010000000010000000100",
		1181 =>	"00000100000001000000010000001000",
		1182 =>	"00001110000001000000010000000100",
		1183 =>	"00000100000001000000001100000011",
		1184 =>	"00000011000011100000111000000100",
		1185 =>	"00001000000001000000010000001000",
		1186 =>	"00001110000001000000010000001110",
		1187 =>	"00001110000011100000001100000011",
		1188 =>	"00000011000010000000010000000100",
		1189 =>	"00001000000001000000010000001000",
		1190 =>	"00001110000010000000010000001110",
		1191 =>	"00000100000001000000001100000011",
		1192 =>	"00000011000011100000111000000100",
		1193 =>	"00001000000010000000010000001000",
		1194 =>	"00001110000010000000111000001110",
		1195 =>	"00001110000011100000001100000011",
		1196 =>	"00000011000010000000010000000100",
		1197 =>	"00001000000010000000100000001000",
		1198 =>	"00001000000010000000111000001110",
		1199 =>	"00000100000001000000001100000011",
		1200 =>	"00000011000011100000111000000100",
		1201 =>	"00001000000001000000010000001110",
		1202 =>	"00000100000001000000111000001110",
		1203 =>	"00001110000011100000001100000011",
		1204 =>	"00000011000010000000010000000100",
		1205 =>	"00001000000001000000111000001110",
		1206 =>	"00001000000001000000111000001110",
		1207 =>	"00000100000001000000001100000011",
		1208 =>	"00000011000011100000111000000100",
		1209 =>	"00001000000001000000111000001000",
		1210 =>	"00001000000001000000111000001110",
		1211 =>	"00001110000011100000001100000011",
		1212 =>	"00000011000010000000010000000100",
		1213 =>	"00001000000001000000010000000100",
		1214 =>	"00000100000001000000111000001110",
		1215 =>	"00000100000001000000001100000011",
		1216 =>	"00000011000011100000111000000100",
		1217 =>	"00001000000001000000010000000100",
		1218 =>	"00000100000001000000111000001110",
		1219 =>	"00001110000011100000001100000011",
		1220 =>	"00000011000010000000010000000100",
		1221 =>	"00000100000011100000111000001110",
		1222 =>	"00001110000011100000010000001110",
		1223 =>	"00000100000001000000001100000011",
		1224 =>	"00000011000011100000111000000100",
		1225 =>	"00001110000011100000111000001110",
		1226 =>	"00001110000011100000111000000100",
		1227 =>	"00001110000011100000001100000011",
		1228 =>	"00000011000010000000010000000100",
		1229 =>	"00000011000000110000001100000100",
		1230 =>	"00000011000000110000001100001110",
		1231 =>	"00000100000001000000001100000011",
		1232 =>	"00000011000000110000001100000011", -- IMG_16x16_EXPLOSION
		1233 =>	"00001111000000110000111100000011",
		1234 =>	"00000011000000110000001100001111",
		1235 =>	"00000011000000110000111100000011",
		1236 =>	"00000011000010000000001100000011",
		1237 =>	"00000011000010000000001100000011",
		1238 =>	"00001000000000110000111100000011",
		1239 =>	"00000011000010000000111100000011",
		1240 =>	"00000011000011110000111100001000",
		1241 =>	"00001000000000110000001100001000",
		1242 =>	"00001000000000110000001100000011",
		1243 =>	"00001000000011110000001100000011",
		1244 =>	"00000011000000110000111100001111",
		1245 =>	"00001000000011110000111100001000",
		1246 =>	"00001111000011110000001100001000",
		1247 =>	"00001000000011110000001100000011",
		1248 =>	"00000011000000110000001100001111",
		1249 =>	"00010000000010000000100000001000",
		1250 =>	"00001000000011110000100000001000",
		1251 =>	"00001111000011110000001100001111",
		1252 =>	"00000011000010000000001100001111",
		1253 =>	"00001000000010000001000000001000",
		1254 =>	"00000011000010000000100000010000",
		1255 =>	"00001111000000110000001100000011",
		1256 =>	"00000011000000110000111100001000",
		1257 =>	"00001000000100000000111100010000",
		1258 =>	"00010000000000110001000000001111",
		1259 =>	"00001000000011110000001100000011",
		1260 =>	"00001000000010000000100000001000",
		1261 =>	"00000011000010000001000000000011",
		1262 =>	"00000011000100000000100000001000",
		1263 =>	"00001000000010000000100000001000",
		1264 =>	"00000011000011110000111100001111",
		1265 =>	"00001000000010000000111100010000",
		1266 =>	"00000011000100000000100000001111",
		1267 =>	"00001111000011110000001100000011",
		1268 =>	"00000011000000110000001100001111",
		1269 =>	"00001111000011110000001100001000",
		1270 =>	"00010000000000110000111100001111",
		1271 =>	"00001000000010000000001100000011",
		1272 =>	"00000011000010000000111100001111",
		1273 =>	"00001000000010000000111100001000",
		1274 =>	"00000011000010000001000000001000",
		1275 =>	"00001111000011110000100000000011",
		1276 =>	"00000011000000110000100000001000",
		1277 =>	"00001000000100000000100000001111",
		1278 =>	"00001000000011110000100000001000",
		1279 =>	"00000011000000110000001100000011",
		1280 =>	"00000011000011110000100000001111",
		1281 =>	"00001111000010000000111100001000",
		1282 =>	"00001000000011110000111100001000",
		1283 =>	"00001000000000110000111100000011",
		1284 =>	"00000011000010000000111100000011",
		1285 =>	"00000011000011110000001100001111",
		1286 =>	"00001000000011110000001100001111",
		1287 =>	"00001111000010000000001100000011",
		1288 =>	"00001000000011110000001100000011",
		1289 =>	"00001111000000110000001100000011",
		1290 =>	"00001000000000110000001100000011",
		1291 =>	"00000011000011110000100000000011",
		1292 =>	"00000011000000110000001100000011",
		1293 =>	"00000011000000110000001100000011",
		1294 =>	"00001000000000110000111100000011",
		1295 =>	"00000011000000110000111100000011",
		1296 =>	"00000011000000110000000100000001", -- IMG_16x16_FLAG
		1297 =>	"00000001000000010000000100000001",
		1298 =>	"00000001000000010000000100000001",
		1299 =>	"00000001000000010000000100000001",
		1300 =>	"00000011000000110000001000000010",
		1301 =>	"00000001000000010000000100000001",
		1302 =>	"00000001000000010000000100000001",
		1303 =>	"00000001000000010000000100000001",
		1304 =>	"00000011000000110000001000000010",
		1305 =>	"00000010000000100000000100000001",
		1306 =>	"00000001000000010000000100000001",
		1307 =>	"00000001000000010000000100000001",
		1308 =>	"00000011000000110000001000000010",
		1309 =>	"00000010000000100000001000000010",
		1310 =>	"00000001000000010000000100000001",
		1311 =>	"00000001000000010000000100000001",
		1312 =>	"00000011000000110000001000000010",
		1313 =>	"00000010000000100000001000000010",
		1314 =>	"00000010000000100000000100000001",
		1315 =>	"00000001000000010000000100000001",
		1316 =>	"00000011000000110000001000000010",
		1317 =>	"00000010000000100000001000000010",
		1318 =>	"00000010000000100000001000000010",
		1319 =>	"00000001000000010000000100000001",
		1320 =>	"00000011000000110000001000000010",
		1321 =>	"00000010000000100000001000000010",
		1322 =>	"00000010000000100000001000000010",
		1323 =>	"00000010000000100000000100000001",
		1324 =>	"00000011000000110000001000000010",
		1325 =>	"00000010000000100000001000000010",
		1326 =>	"00000010000000100000001000000010",
		1327 =>	"00000010000000100000001000000010",
		1328 =>	"00000011000000110000001000000010",
		1329 =>	"00000010000000100000001000000010",
		1330 =>	"00000010000000100000001000000010",
		1331 =>	"00000010000000100000001000000010",
		1332 =>	"00000011000000110000000100000001",
		1333 =>	"00000001000000010000000100000001",
		1334 =>	"00000001000000010000000100000001",
		1335 =>	"00000001000000010000000100000001",
		1336 =>	"00000011000000110000000100000001",
		1337 =>	"00000001000000010000000100000001",
		1338 =>	"00000001000000010000000100000001",
		1339 =>	"00000001000000010000000100000001",
		1340 =>	"00000011000000110000000100000001",
		1341 =>	"00000001000000010000000100000001",
		1342 =>	"00000001000000010000000100000001",
		1343 =>	"00000001000000010000000100000001",
		1344 =>	"00000011000000110000000100000001",
		1345 =>	"00000001000000010000000100000001",
		1346 =>	"00000001000000010000000100000001",
		1347 =>	"00000001000000010000000100000001",
		1348 =>	"00000011000000110000000100000001",
		1349 =>	"00000001000000010000000100000001",
		1350 =>	"00000001000000010000000100000001",
		1351 =>	"00000001000000010000000100000001",
		1352 =>	"00000011000000110000000100000001",
		1353 =>	"00000001000000010000000100000001",
		1354 =>	"00000001000000010000000100000001",
		1355 =>	"00000001000000010000000100000001",
		1356 =>	"00000001000000010000000100000001",
		1357 =>	"00000001000000010000000100000001",
		1358 =>	"00000001000000010000000100000001",
		1359 =>	"00000001000000010000000100000001",
		1360 =>	"00000011000000110000001100000011", -- IMG_16x16_MAIN_TANK
		1361 =>	"00000011000000110000001100000011",
		1362 =>	"00000011000000110000001100000011",
		1363 =>	"00000011000000110000001100000011",
		1364 =>	"00000011000000110000001100000011",
		1365 =>	"00000011000000110000001100000011",
		1366 =>	"00000011000000110000001100000011",
		1367 =>	"00000011000000110000001100000011",
		1368 =>	"00000011000000110000001100000011",
		1369 =>	"00000011000000110000001100010001",
		1370 =>	"00000011000000110000001100000011",
		1371 =>	"00000011000000110000001100000011",
		1372 =>	"00000011000000110000001100000011",
		1373 =>	"00000011000000110000001100010001",
		1374 =>	"00000011000000110000001100000011",
		1375 =>	"00000011000000110000001100000011",
		1376 =>	"00000011000100010001001000010010",
		1377 =>	"00000011000000110000001100010001",
		1378 =>	"00000011000000110000001100010001",
		1379 =>	"00010010000100100000001100000011",
		1380 =>	"00000011000100110001001100010001",
		1381 =>	"00000011000000110000001100010001",
		1382 =>	"00000011000000110000001100010011",
		1383 =>	"00010011000100110000001100000011",
		1384 =>	"00000011000100010001001000010001",
		1385 =>	"00000011000100010001001000010001",
		1386 =>	"00010011000100110000001100010011",
		1387 =>	"00010010000100100000001100000011",
		1388 =>	"00000011000100110001001100010001",
		1389 =>	"00010001000100010001001000010010",
		1390 =>	"00010010000100100001001100010011",
		1391 =>	"00010011000100110000001100000011",
		1392 =>	"00000011000100010001001000010001",
		1393 =>	"00010001000100100001000100010001",
		1394 =>	"00010010000100100001001000010011",
		1395 =>	"00010010000100100000001100000011",
		1396 =>	"00000011000100110001001100010001",
		1397 =>	"00010001000100100001000100010010",
		1398 =>	"00010011000100100001001000010011",
		1399 =>	"00010011000100110000001100000011",
		1400 =>	"00000011000100010001001000010001",
		1401 =>	"00010001000100100001000100010010",
		1402 =>	"00010011000100100001001000010011",
		1403 =>	"00010010000100100000001100000011",
		1404 =>	"00000011000100110001001100010001",
		1405 =>	"00010001000100010001001000010011",
		1406 =>	"00010011000100100001001000010011",
		1407 =>	"00010011000100110000001100000011",
		1408 =>	"00000011000100010001001000010001",
		1409 =>	"00010011000100010001000100010010",
		1410 =>	"00010010000100100001001100010011",
		1411 =>	"00010010000100100000001100000011",
		1412 =>	"00000011000100110001001100010001",
		1413 =>	"00000011000100110001001100010011",
		1414 =>	"00010011000100110000001100010011",
		1415 =>	"00010011000100110000001100000011",
		1416 =>	"00000011000100010001001000010010",
		1417 =>	"00000011000000110000001100000011",
		1418 =>	"00000011000000110000001100010011",
		1419 =>	"00010010000100100000001100000011",
		1420 =>	"00000011000000110000001100000011",
		1421 =>	"00000011000000110000001100000011",
		1422 =>	"00000011000000110000001100000011",
		1423 =>	"00000011000000110000001100000011",


--			***** MAP *****


		1424 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 256
		1425 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 272
		1426 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 288
		1427 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 304
		1428 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 320
		1429 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 336
		1430 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 352
		1431 =>	"00000000000000000000000101100000", -- z: 1 rot: 0 ptr: 368
		1432 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1433 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1434 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1435 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1436 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1437 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1438 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1439 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1440 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1441 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1442 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1443 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1444 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1445 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1446 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1447 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1448 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1449 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1450 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1451 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1452 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1453 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1454 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1455 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1456 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1457 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1458 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1459 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1460 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1461 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1462 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1463 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1464 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1465 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1466 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1467 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1468 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1469 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1470 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1471 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1472 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1473 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1474 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1475 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1476 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1477 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1478 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1479 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1480 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1481 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1482 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1483 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1484 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1485 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1486 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1487 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1488 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1489 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1490 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1491 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1492 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1493 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1494 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1495 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1496 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1497 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1498 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1499 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1500 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1501 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1502 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1503 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1504 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1505 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1506 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1507 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1508 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1509 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1510 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1511 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1512 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1513 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1514 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1515 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1516 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1517 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1518 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1519 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1520 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1521 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1522 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1523 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1524 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1525 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1526 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1527 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1528 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1529 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1530 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1531 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1532 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1533 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1534 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1535 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1536 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1537 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1538 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1539 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1540 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1541 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1542 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1543 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1544 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1545 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1546 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1547 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1548 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1549 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1550 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1551 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1552 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1553 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1554 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1555 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1556 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1557 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1558 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1559 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1560 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1561 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1562 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1563 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1564 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1565 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1566 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1567 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1568 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1569 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1570 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1571 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1572 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1573 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1574 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1575 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1576 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1577 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1578 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1579 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1580 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1581 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1582 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1583 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1584 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1585 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1586 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1587 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1588 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1589 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1590 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1591 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1592 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1593 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1594 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1595 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1596 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1597 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1598 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1599 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1600 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1601 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1602 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1603 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1604 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1605 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1606 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1607 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1608 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1609 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1610 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1611 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1612 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1613 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1614 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1615 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1616 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1617 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1618 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1619 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1620 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1621 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1622 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1623 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1624 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1625 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1626 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1627 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1628 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1629 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1630 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1631 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1632 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1633 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1634 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1635 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1636 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1637 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1638 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1639 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1640 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1641 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1642 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1643 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1644 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1645 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1646 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1647 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1648 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1649 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1650 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1651 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1652 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1653 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1654 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1655 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1656 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1657 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1658 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1659 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1660 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1661 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1662 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1663 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1664 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1665 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1666 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1667 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1668 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1669 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1670 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1671 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1672 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1673 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1674 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1675 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1676 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1677 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1678 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1679 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1680 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1681 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1682 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1683 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1684 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1685 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1686 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1687 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1688 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1689 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1690 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1691 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1692 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1693 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1694 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1695 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1696 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1697 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1698 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1699 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1700 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1701 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1702 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1703 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1704 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1705 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1706 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1707 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1708 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1709 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1710 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1711 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1712 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1713 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1714 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1715 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1716 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1717 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1718 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1719 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1720 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1721 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1722 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1723 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1724 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1725 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1726 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1727 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1728 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1729 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1730 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1731 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1732 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1733 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1734 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1735 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1736 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1737 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1738 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1739 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1740 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1741 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1742 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1743 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1744 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1745 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1746 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1747 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1748 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1749 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1750 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1751 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1752 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1753 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1754 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1755 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1756 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1757 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1758 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1759 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1760 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1761 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1762 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1763 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1764 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1765 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1766 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1767 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1768 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1769 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1770 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1771 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1772 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1773 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1774 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1775 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1776 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1777 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1778 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1779 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1780 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1781 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1782 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1783 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1784 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1785 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1786 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1787 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1788 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1789 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1790 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1791 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1792 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1793 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1794 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1795 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1796 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1797 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1798 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1799 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1800 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1801 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1802 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1803 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1804 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1805 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1806 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1807 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1808 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1809 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1810 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1811 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1812 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1813 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1814 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1815 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1816 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1817 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1818 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1819 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1820 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1821 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1822 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1823 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1824 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1825 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1826 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1827 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1828 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1829 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1830 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1831 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1832 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1833 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1834 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1835 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1836 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1837 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1838 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1839 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1840 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1841 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1842 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1843 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1844 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1845 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1846 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1847 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1848 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1849 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1850 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1851 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1852 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1853 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1854 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1855 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1856 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1857 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1858 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1859 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1860 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1861 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1862 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1863 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1864 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1865 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1866 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1867 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1868 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1869 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1870 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1871 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1872 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1873 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1874 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1875 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1876 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1877 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1878 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1879 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1880 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1881 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1882 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1883 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1884 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1885 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1886 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1887 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1888 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1889 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1890 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1891 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1892 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1893 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1894 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1895 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1896 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1897 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1898 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1899 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1900 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1901 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1902 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1903 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1904 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1905 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1906 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1907 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1908 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1909 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1910 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1911 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1912 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1913 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1914 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1915 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1916 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1917 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1918 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1919 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1920 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1921 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1922 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1923 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1924 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1925 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1926 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1927 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1928 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1929 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1930 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1931 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1932 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1933 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1934 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1935 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1936 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1937 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1938 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1939 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1940 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1941 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1942 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1943 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1944 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1945 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1946 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1947 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1948 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1949 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1950 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1951 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1952 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1953 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1954 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1955 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1956 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1957 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1958 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1959 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1960 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1961 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1962 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1963 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1964 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1965 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1966 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1967 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1968 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1969 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1970 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1971 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1972 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1973 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1974 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1975 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1976 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1977 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1978 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1979 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1980 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1981 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1982 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1983 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1984 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1985 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1986 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1987 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1988 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1989 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1990 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1991 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1992 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1993 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1994 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1995 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1996 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1997 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1998 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		1999 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2000 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2001 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2002 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2003 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2004 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2005 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2006 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2007 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2008 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2009 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2010 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2011 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2012 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2013 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2014 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2015 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2016 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2017 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2018 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2019 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2020 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2021 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2022 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2023 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2024 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2025 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2026 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2027 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2028 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2029 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2030 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2031 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2032 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2033 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2034 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2035 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2036 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2037 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2038 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2039 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2040 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2041 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2042 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2043 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2044 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2045 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2046 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2047 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2048 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2049 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2050 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2051 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2052 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2053 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2054 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2055 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2056 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2057 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2058 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2059 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2060 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2061 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2062 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2063 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2064 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2065 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2066 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2067 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2068 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2069 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2070 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2071 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2072 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2073 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2074 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2075 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2076 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2077 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2078 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2079 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2080 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2081 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2082 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2083 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2084 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2085 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2086 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2087 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2088 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2089 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2090 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2091 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2092 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2093 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2094 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2095 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2096 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2097 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2098 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2099 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2100 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2101 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2102 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2103 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2104 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2105 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2106 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2107 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2108 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2109 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2110 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2111 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2112 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2113 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2114 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2115 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2116 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2117 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2118 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2119 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2120 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2121 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2122 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2123 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2124 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2125 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2126 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2127 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2128 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2129 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2130 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2131 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2132 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2133 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2134 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2135 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2136 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2137 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2138 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2139 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2140 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2141 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2142 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2143 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2144 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2145 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2146 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2147 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2148 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2149 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2150 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2151 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2152 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2153 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2154 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2155 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2156 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2157 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2158 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2159 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2160 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2161 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2162 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2163 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2164 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2165 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2166 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2167 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2168 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2169 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2170 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2171 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2172 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2173 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2174 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2175 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2176 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2177 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2178 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2179 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2180 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2181 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2182 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2183 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2184 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2185 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2186 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2187 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2188 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2189 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2190 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2191 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2192 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2193 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2194 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2195 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2196 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2197 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2198 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2199 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2200 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2201 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2202 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2203 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2204 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2205 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2206 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2207 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2208 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2209 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2210 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2211 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2212 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2213 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2214 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2215 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2216 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2217 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2218 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2219 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2220 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2221 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2222 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2223 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2224 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2225 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2226 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2227 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2228 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2229 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2230 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2231 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2232 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2233 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2234 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2235 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2236 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2237 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2238 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2239 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2240 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2241 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2242 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2243 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2244 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2245 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2246 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2247 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2248 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2249 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2250 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2251 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2252 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2253 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2254 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2255 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2256 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2257 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2258 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2259 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2260 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2261 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2262 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2263 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2264 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2265 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2266 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2267 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2268 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2269 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2270 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2271 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2272 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2273 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2274 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2275 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2276 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2277 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2278 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2279 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2280 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2281 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2282 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2283 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2284 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2285 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2286 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2287 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2288 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2289 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2290 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2291 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2292 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2293 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2294 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2295 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2296 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2297 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2298 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2299 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2300 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2301 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2302 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2303 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2304 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2305 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2306 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2307 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2308 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2309 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2310 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2311 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2312 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2313 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2314 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2315 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2316 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2317 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2318 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2319 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2320 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2321 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2322 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2323 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2324 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2325 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2326 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2327 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2328 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2329 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2330 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2331 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2332 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2333 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2334 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2335 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2336 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2337 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2338 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2339 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2340 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2341 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2342 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2343 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2344 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2345 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2346 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2347 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2348 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2349 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2350 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2351 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2352 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2353 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2354 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2355 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2356 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2357 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2358 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2359 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2360 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2361 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2362 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2363 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2364 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2365 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2366 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2367 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2368 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2369 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2370 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2371 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2372 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2373 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2374 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2375 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2376 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2377 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2378 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2379 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2380 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2381 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2382 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2383 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2384 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2385 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2386 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2387 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2388 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2389 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2390 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2391 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2392 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2393 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2394 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2395 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2396 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2397 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2398 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2399 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2400 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2401 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2402 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2403 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2404 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2405 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2406 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2407 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2408 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2409 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2410 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2411 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2412 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2413 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2414 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2415 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2416 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2417 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2418 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2419 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2420 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2421 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2422 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2423 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2424 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2425 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2426 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2427 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2428 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2429 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2430 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2431 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2432 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2433 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2434 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2435 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2436 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2437 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2438 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2439 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2440 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2441 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2442 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2443 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2444 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2445 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2446 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2447 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2448 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2449 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2450 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2451 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2452 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2453 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2454 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2455 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2456 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2457 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2458 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2459 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2460 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2461 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2462 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2463 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2464 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2465 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2466 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2467 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2468 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2469 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2470 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2471 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2472 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2473 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2474 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2475 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2476 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2477 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2478 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2479 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2480 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2481 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2482 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2483 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2484 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2485 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2486 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2487 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2488 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2489 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2490 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2491 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2492 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2493 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2494 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2495 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2496 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2497 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2498 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2499 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2500 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2501 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2502 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2503 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2504 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2505 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2506 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2507 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2508 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2509 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2510 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2511 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2512 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2513 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2514 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2515 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2516 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2517 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2518 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2519 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2520 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2521 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2522 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2523 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2524 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2525 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2526 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2527 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2528 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2529 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2530 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2531 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2532 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2533 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2534 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2535 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2536 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2537 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2538 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2539 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2540 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2541 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2542 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2543 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2544 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2545 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2546 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2547 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2548 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2549 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2550 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2551 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2552 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2553 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2554 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2555 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2556 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2557 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2558 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2559 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2560 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2561 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2562 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2563 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2564 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2565 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2566 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2567 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2568 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2569 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2570 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2571 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2572 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2573 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2574 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2575 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2576 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2577 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2578 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2579 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2580 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2581 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2582 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2583 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2584 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2585 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2586 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2587 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2588 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2589 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2590 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2591 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2592 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2593 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2594 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2595 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2596 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2597 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2598 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2599 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2600 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2601 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2602 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2603 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2604 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2605 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2606 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2607 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2608 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2609 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2610 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2611 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2612 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2613 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2614 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2615 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2616 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2617 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2618 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2619 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2620 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2621 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2622 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2623 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2624 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2625 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2626 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2627 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2628 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2629 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2630 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2631 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2632 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2633 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2634 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2635 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2636 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2637 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2638 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2639 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2640 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2641 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2642 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2643 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2644 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2645 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2646 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2647 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2648 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2649 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2650 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2651 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2652 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2653 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2654 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2655 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2656 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2657 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2658 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2659 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2660 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2661 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2662 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2663 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2664 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2665 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2666 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2667 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2668 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2669 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2670 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2671 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2672 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2673 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2674 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2675 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2676 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2677 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2678 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2679 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2680 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2681 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2682 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2683 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2684 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2685 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2686 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2687 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2688 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2689 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2690 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2691 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2692 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2693 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2694 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2695 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2696 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2697 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2698 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2699 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2700 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2701 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2702 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2703 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2704 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2705 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2706 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2707 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2708 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2709 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2710 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2711 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2712 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2713 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2714 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2715 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2716 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2717 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2718 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2719 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2720 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2721 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2722 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2723 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2724 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2725 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2726 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2727 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2728 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2729 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2730 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2731 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2732 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2733 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2734 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2735 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2736 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2737 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2738 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2739 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2740 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2741 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2742 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2743 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2744 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2745 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2746 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2747 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2748 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2749 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2750 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2751 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2752 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2753 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2754 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2755 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2756 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2757 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2758 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2759 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2760 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2761 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2762 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2763 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2764 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2765 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2766 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2767 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2768 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2769 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2770 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2771 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2772 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2773 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2774 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2775 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2776 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2777 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2778 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2779 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2780 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2781 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2782 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2783 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2784 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2785 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2786 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2787 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2788 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2789 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2790 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2791 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2792 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2793 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2794 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2795 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2796 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2797 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2798 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2799 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2800 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2801 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2802 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2803 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2804 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2805 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2806 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2807 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2808 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2809 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2810 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2811 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2812 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2813 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2814 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2815 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2816 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2817 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2818 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2819 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2820 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2821 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2822 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2823 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2824 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2825 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2826 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2827 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2828 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2829 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2830 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2831 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2832 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2833 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2834 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2835 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2836 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2837 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2838 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2839 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2840 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2841 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2842 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2843 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2844 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2845 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2846 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2847 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2848 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2849 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2850 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2851 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2852 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2853 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2854 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2855 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2856 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2857 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2858 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2859 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2860 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2861 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2862 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2863 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2864 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2865 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2866 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2867 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2868 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2869 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2870 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2871 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2872 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2873 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2874 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2875 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2876 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2877 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2878 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2879 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2880 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2881 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2882 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2883 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2884 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2885 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2886 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2887 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2888 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2889 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2890 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2891 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2892 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2893 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2894 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2895 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2896 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2897 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2898 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2899 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2900 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2901 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2902 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2903 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2904 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2905 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2906 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2907 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2908 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2909 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2910 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2911 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2912 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2913 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2914 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2915 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2916 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2917 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2918 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2919 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2920 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2921 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2922 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2923 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2924 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2925 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2926 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2927 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2928 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2929 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2930 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2931 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2932 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2933 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2934 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2935 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2936 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2937 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2938 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2939 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2940 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2941 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2942 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2943 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2944 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2945 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2946 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2947 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2948 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2949 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2950 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2951 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2952 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2953 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2954 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2955 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2956 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2957 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2958 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2959 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2960 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2961 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2962 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2963 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2964 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2965 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2966 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2967 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2968 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2969 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2970 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2971 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2972 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2973 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2974 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2975 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2976 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2977 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2978 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2979 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2980 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2981 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2982 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2983 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2984 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2985 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2986 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2987 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2988 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2989 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2990 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2991 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2992 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2993 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2994 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2995 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2996 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2997 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2998 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		2999 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3000 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3001 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3002 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3003 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3004 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3005 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3006 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3007 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3008 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3009 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3010 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3011 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3012 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3013 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3014 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3015 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3016 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3017 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3018 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3019 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3020 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3021 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3022 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3023 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3024 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3025 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3026 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3027 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3028 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3029 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3030 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3031 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3032 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3033 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3034 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3035 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3036 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3037 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3038 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3039 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3040 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3041 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3042 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3043 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3044 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3045 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3046 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3047 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3048 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3049 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3050 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3051 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3052 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3053 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3054 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3055 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3056 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3057 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3058 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3059 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3060 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3061 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3062 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3063 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3064 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3065 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3066 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3067 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3068 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3069 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3070 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3071 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3072 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3073 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3074 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3075 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3076 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3077 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3078 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3079 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3080 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3081 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3082 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3083 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3084 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3085 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3086 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3087 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3088 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3089 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3090 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3091 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3092 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3093 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3094 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3095 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3096 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3097 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3098 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3099 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3100 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3101 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3102 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3103 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3104 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3105 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3106 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3107 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3108 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3109 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3110 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3111 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3112 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3113 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3114 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3115 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3116 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3117 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3118 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3119 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3120 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3121 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3122 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3123 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3124 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3125 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3126 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3127 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3128 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3129 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3130 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3131 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3132 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3133 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3134 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3135 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3136 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3137 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3138 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3139 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3140 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3141 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3142 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3143 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3144 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3145 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3146 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3147 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3148 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3149 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3150 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3151 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3152 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3153 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3154 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3155 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3156 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3157 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3158 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3159 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3160 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3161 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3162 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3163 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3164 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3165 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3166 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3167 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3168 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3169 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3170 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3171 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3172 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3173 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3174 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3175 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3176 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3177 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3178 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3179 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3180 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3181 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3182 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3183 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3184 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3185 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3186 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3187 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3188 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3189 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3190 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3191 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3192 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3193 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3194 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3195 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3196 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3197 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3198 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3199 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3200 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3201 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3202 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3203 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3204 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3205 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3206 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3207 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3208 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3209 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3210 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3211 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3212 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3213 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3214 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3215 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3216 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3217 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3218 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3219 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3220 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3221 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3222 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3223 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3224 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3225 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3226 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3227 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3228 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3229 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3230 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3231 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3232 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3233 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3234 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3235 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3236 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3237 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3238 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3239 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3240 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3241 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3242 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3243 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3244 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3245 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3246 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3247 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3248 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3249 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3250 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3251 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3252 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3253 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3254 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3255 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3256 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3257 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3258 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3259 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3260 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3261 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3262 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3263 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3264 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3265 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3266 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3267 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3268 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3269 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3270 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3271 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3272 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3273 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3274 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3275 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3276 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3277 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3278 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3279 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3280 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3281 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3282 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3283 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3284 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3285 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3286 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3287 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3288 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3289 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3290 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3291 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3292 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3293 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3294 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3295 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3296 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3297 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3298 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3299 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3300 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3301 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3302 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3303 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3304 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3305 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3306 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3307 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3308 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3309 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3310 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3311 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3312 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3313 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3314 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3315 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3316 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3317 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3318 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3319 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3320 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3321 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3322 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3323 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3324 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3325 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3326 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3327 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3328 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3329 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3330 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3331 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3332 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3333 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3334 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3335 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3336 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3337 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3338 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3339 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3340 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3341 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3342 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3343 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3344 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3345 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3346 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3347 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3348 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3349 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3350 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3351 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3352 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3353 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3354 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3355 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3356 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3357 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3358 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3359 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3360 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3361 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3362 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3363 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3364 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3365 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3366 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3367 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3368 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3369 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3370 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3371 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3372 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3373 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3374 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3375 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3376 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3377 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3378 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3379 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3380 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3381 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3382 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3383 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3384 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3385 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3386 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3387 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3388 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3389 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3390 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3391 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3392 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3393 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3394 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3395 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3396 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3397 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3398 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3399 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3400 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3401 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3402 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3403 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3404 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3405 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3406 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3407 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3408 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3409 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3410 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3411 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3412 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3413 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3414 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3415 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3416 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3417 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3418 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3419 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3420 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3421 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3422 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3423 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3424 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3425 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3426 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3427 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3428 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3429 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3430 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3431 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3432 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3433 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3434 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3435 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3436 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3437 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3438 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3439 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3440 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3441 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3442 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3443 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3444 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3445 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3446 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3447 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3448 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3449 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3450 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3451 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3452 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3453 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3454 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3455 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3456 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3457 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3458 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3459 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3460 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3461 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3462 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3463 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3464 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3465 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3466 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3467 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3468 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3469 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3470 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3471 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3472 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3473 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3474 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3475 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3476 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3477 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3478 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3479 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3480 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3481 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3482 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3483 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3484 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3485 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3486 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3487 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3488 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3489 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3490 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3491 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3492 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3493 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3494 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3495 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3496 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3497 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3498 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3499 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3500 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3501 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3502 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3503 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3504 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3505 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3506 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3507 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3508 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3509 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3510 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3511 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3512 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3513 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3514 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3515 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3516 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3517 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3518 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3519 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3520 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3521 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3522 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3523 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3524 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3525 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3526 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3527 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3528 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3529 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3530 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3531 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3532 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3533 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3534 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3535 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3536 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3537 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3538 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3539 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3540 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3541 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3542 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3543 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3544 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3545 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3546 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3547 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3548 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3549 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3550 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3551 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3552 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3553 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3554 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3555 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3556 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3557 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3558 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3559 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3560 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3561 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3562 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3563 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3564 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3565 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3566 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3567 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3568 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3569 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3570 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3571 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3572 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3573 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3574 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3575 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3576 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3577 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3578 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3579 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3580 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3581 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3582 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3583 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3584 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3585 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3586 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3587 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3588 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3589 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3590 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3591 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3592 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3593 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3594 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3595 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3596 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3597 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3598 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3599 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3600 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3601 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3602 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3603 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3604 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3605 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3606 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3607 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3608 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3609 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3610 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3611 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3612 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3613 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3614 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3615 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3616 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3617 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3618 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3619 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3620 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3621 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3622 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3623 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3624 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3625 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3626 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3627 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3628 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3629 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3630 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3631 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3632 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3633 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3634 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3635 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3636 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3637 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3638 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3639 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3640 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3641 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3642 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3643 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3644 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3645 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3646 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3647 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3648 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3649 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3650 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3651 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3652 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3653 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3654 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3655 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3656 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3657 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3658 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3659 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3660 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3661 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3662 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3663 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3664 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3665 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3666 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3667 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3668 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3669 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3670 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3671 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3672 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3673 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3674 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3675 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3676 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3677 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3678 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3679 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3680 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3681 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3682 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3683 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3684 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3685 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3686 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3687 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3688 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3689 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3690 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3691 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3692 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3693 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3694 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3695 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3696 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3697 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3698 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3699 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3700 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3701 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3702 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3703 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3704 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3705 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3706 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3707 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3708 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3709 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3710 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3711 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3712 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3713 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3714 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3715 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3716 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3717 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3718 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3719 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3720 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3721 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3722 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3723 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3724 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3725 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3726 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3727 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3728 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3729 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3730 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3731 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3732 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3733 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3734 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3735 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3736 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3737 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3738 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3739 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3740 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3741 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3742 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3743 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3744 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3745 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3746 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3747 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3748 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3749 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3750 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3751 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3752 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3753 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3754 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3755 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3756 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3757 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3758 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3759 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3760 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3761 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3762 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3763 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3764 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3765 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3766 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3767 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3768 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3769 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3770 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3771 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3772 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3773 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3774 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3775 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3776 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3777 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3778 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3779 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3780 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3781 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3782 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3783 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3784 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3785 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3786 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3787 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3788 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3789 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3790 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3791 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3792 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3793 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3794 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3795 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3796 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3797 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3798 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3799 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3800 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3801 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3802 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3803 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3804 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3805 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3806 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3807 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3808 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3809 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3810 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3811 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3812 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3813 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3814 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3815 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3816 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3817 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3818 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3819 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3820 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3821 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3822 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3823 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3824 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3825 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3826 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3827 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3828 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3829 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3830 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3831 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3832 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3833 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3834 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3835 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3836 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3837 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3838 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3839 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3840 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3841 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3842 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3843 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3844 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3845 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3846 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3847 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3848 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3849 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3850 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3851 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3852 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3853 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3854 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3855 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3856 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3857 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3858 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3859 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3860 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3861 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3862 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3863 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3864 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3865 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3866 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3867 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3868 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3869 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3870 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3871 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3872 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3873 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3874 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3875 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3876 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3877 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3878 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3879 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3880 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3881 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3882 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3883 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3884 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3885 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3886 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3887 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3888 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3889 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3890 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3891 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3892 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3893 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3894 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3895 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3896 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3897 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3898 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3899 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3900 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3901 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3902 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3903 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3904 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3905 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3906 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3907 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3908 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3909 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3910 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3911 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3912 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3913 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3914 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3915 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3916 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3917 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3918 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3919 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3920 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3921 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3922 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3923 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3924 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3925 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3926 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3927 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3928 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3929 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3930 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3931 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3932 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3933 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3934 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3935 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3936 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3937 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3938 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3939 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3940 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3941 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3942 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3943 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3944 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3945 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3946 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3947 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3948 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3949 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3950 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3951 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3952 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3953 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3954 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3955 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3956 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3957 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3958 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3959 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3960 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3961 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3962 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3963 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3964 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3965 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3966 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3967 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3968 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3969 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3970 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3971 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3972 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3973 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3974 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3975 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3976 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3977 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3978 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3979 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3980 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3981 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3982 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3983 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3984 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3985 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3986 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3987 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3988 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3989 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3990 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3991 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3992 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3993 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3994 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3995 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3996 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3997 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3998 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		3999 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4000 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4001 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4002 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4003 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4004 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4005 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4006 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4007 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4008 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4009 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4010 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4011 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4012 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4013 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4014 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4015 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4016 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4017 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4018 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4019 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4020 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4021 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4022 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4023 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4024 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4025 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4026 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4027 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4028 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4029 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4030 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4031 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4032 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4033 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4034 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4035 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4036 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4037 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4038 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4039 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4040 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4041 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4042 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4043 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4044 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4045 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4046 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4047 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4048 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4049 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4050 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4051 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4052 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4053 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4054 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4055 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4056 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4057 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4058 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4059 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4060 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4061 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4062 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4063 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4064 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4065 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4066 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4067 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4068 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4069 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4070 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4071 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4072 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4073 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4074 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4075 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4076 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4077 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4078 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4079 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4080 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4081 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4082 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4083 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4084 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4085 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4086 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4087 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4088 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4089 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4090 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4091 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4092 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4093 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4094 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4095 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4096 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4097 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4098 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4099 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4100 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4101 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4102 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4103 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4104 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4105 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4106 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4107 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4108 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4109 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4110 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4111 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4112 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4113 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4114 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4115 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4116 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4117 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4118 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4119 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4120 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4121 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4122 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4123 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4124 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4125 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4126 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4127 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4128 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4129 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4130 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4131 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4132 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4133 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4134 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4135 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4136 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4137 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4138 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4139 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4140 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4141 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4142 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4143 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4144 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4145 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4146 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4147 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4148 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4149 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4150 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4151 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4152 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4153 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4154 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4155 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4156 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4157 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4158 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4159 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4160 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4161 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4162 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4163 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4164 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4165 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4166 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4167 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4168 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4169 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4170 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4171 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4172 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4173 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4174 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4175 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4176 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4177 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4178 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4179 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4180 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4181 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4182 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4183 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4184 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4185 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4186 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4187 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4188 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4189 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4190 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4191 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4192 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4193 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4194 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4195 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4196 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4197 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4198 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4199 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4200 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4201 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4202 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4203 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4204 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4205 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4206 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4207 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4208 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4209 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4210 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4211 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4212 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4213 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4214 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4215 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4216 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4217 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4218 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4219 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4220 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4221 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4222 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4223 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4224 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4225 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4226 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4227 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4228 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4229 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4230 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4231 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4232 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4233 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4234 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4235 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4236 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4237 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4238 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4239 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4240 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4241 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4242 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4243 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4244 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4245 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4246 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4247 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4248 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4249 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4250 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4251 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4252 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4253 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4254 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4255 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4256 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4257 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4258 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4259 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4260 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4261 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4262 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4263 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4264 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4265 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4266 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4267 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4268 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4269 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4270 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4271 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4272 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4273 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4274 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4275 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4276 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4277 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4278 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4279 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4280 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4281 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4282 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4283 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4284 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4285 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4286 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4287 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4288 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4289 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4290 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4291 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4292 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4293 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4294 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4295 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4296 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4297 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4298 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4299 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4300 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4301 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4302 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4303 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4304 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4305 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4306 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4307 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4308 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4309 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4310 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4311 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4312 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4313 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4314 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4315 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4316 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4317 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4318 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4319 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4320 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4321 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4322 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4323 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4324 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4325 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4326 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4327 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4328 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4329 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4330 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4331 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4332 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4333 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4334 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4335 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4336 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4337 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4338 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4339 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4340 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4341 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4342 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4343 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4344 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4345 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4346 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4347 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4348 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4349 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4350 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4351 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4352 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4353 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4354 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4355 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4356 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4357 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4358 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4359 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4360 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4361 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4362 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4363 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4364 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4365 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4366 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4367 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4368 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4369 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4370 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4371 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4372 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4373 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4374 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4375 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4376 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4377 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4378 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4379 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4380 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4381 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4382 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4383 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4384 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4385 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4386 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4387 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4388 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4389 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4390 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4391 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4392 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4393 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4394 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4395 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4396 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4397 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4398 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4399 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4400 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4401 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4402 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4403 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4404 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4405 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4406 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4407 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4408 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4409 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4410 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4411 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4412 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4413 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4414 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4415 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4416 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4417 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4418 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4419 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4420 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4421 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4422 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4423 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4424 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4425 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4426 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4427 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4428 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4429 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4430 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4431 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4432 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4433 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4434 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4435 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4436 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4437 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4438 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4439 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4440 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4441 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4442 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4443 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4444 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4445 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4446 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4447 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4448 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4449 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4450 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4451 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4452 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4453 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4454 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4455 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4456 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4457 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4458 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4459 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4460 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4461 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4462 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4463 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4464 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4465 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4466 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4467 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4468 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4469 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4470 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4471 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4472 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4473 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4474 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4475 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4476 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4477 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4478 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4479 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4480 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4481 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4482 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4483 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4484 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4485 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4486 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4487 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4488 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4489 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4490 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4491 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4492 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4493 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4494 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4495 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4496 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4497 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4498 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4499 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4500 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4501 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4502 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4503 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4504 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4505 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4506 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4507 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4508 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4509 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4510 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4511 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4512 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4513 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4514 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4515 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4516 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4517 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4518 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4519 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4520 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4521 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4522 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4523 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4524 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4525 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4526 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4527 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4528 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4529 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4530 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4531 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4532 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4533 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4534 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4535 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4536 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4537 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4538 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4539 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4540 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4541 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4542 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4543 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4544 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4545 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4546 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4547 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4548 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4549 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4550 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4551 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4552 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4553 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4554 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4555 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4556 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4557 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4558 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4559 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4560 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4561 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4562 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4563 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4564 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4565 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4566 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4567 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4568 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4569 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4570 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4571 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4572 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4573 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4574 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4575 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4576 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4577 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4578 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4579 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4580 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4581 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4582 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4583 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4584 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4585 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4586 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4587 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4588 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4589 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4590 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4591 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4592 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4593 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4594 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4595 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4596 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4597 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4598 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4599 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4600 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4601 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4602 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4603 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4604 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4605 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4606 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4607 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4608 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4609 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4610 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4611 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4612 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4613 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4614 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4615 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4616 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4617 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4618 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4619 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4620 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4621 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4622 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4623 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4624 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4625 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4626 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4627 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4628 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4629 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4630 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4631 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4632 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4633 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4634 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4635 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4636 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4637 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4638 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4639 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4640 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4641 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4642 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4643 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4644 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4645 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4646 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4647 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4648 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4649 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4650 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4651 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4652 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4653 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4654 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4655 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4656 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4657 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4658 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4659 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4660 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4661 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4662 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4663 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4664 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4665 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4666 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4667 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4668 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4669 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4670 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4671 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4672 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4673 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4674 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4675 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4676 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4677 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4678 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4679 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4680 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4681 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4682 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4683 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4684 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4685 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4686 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4687 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4688 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4689 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4690 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4691 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4692 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4693 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4694 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4695 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4696 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4697 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4698 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4699 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4700 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4701 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4702 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4703 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4704 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4705 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4706 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4707 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4708 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4709 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4710 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4711 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4712 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4713 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4714 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4715 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4716 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4717 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4718 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4719 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4720 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4721 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4722 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4723 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4724 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4725 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4726 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4727 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4728 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4729 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4730 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4731 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4732 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4733 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4734 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4735 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4736 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4737 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4738 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4739 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4740 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4741 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4742 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4743 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4744 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4745 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4746 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4747 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4748 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4749 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4750 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4751 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4752 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4753 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4754 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4755 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4756 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4757 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4758 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4759 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4760 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4761 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4762 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4763 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4764 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4765 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4766 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4767 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4768 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4769 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4770 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4771 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4772 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4773 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4774 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4775 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4776 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4777 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4778 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4779 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4780 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4781 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4782 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4783 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4784 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4785 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4786 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4787 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4788 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4789 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4790 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4791 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4792 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4793 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4794 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4795 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4796 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4797 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4798 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4799 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4800 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4801 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4802 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4803 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4804 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4805 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4806 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4807 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4808 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4809 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4810 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4811 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4812 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4813 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4814 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4815 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4816 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4817 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4818 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4819 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4820 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4821 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4822 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4823 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4824 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4825 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4826 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4827 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4828 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4829 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4830 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4831 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4832 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4833 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4834 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4835 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4836 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4837 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4838 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4839 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4840 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4841 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4842 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4843 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4844 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4845 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4846 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4847 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4848 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4849 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4850 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4851 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4852 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4853 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4854 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4855 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4856 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4857 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4858 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4859 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4860 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4861 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4862 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4863 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4864 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4865 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4866 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4867 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4868 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4869 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4870 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4871 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4872 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4873 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4874 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4875 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4876 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4877 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4878 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4879 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4880 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4881 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4882 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4883 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4884 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4885 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4886 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4887 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4888 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4889 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4890 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4891 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4892 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4893 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4894 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4895 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4896 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4897 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4898 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4899 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4900 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4901 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4902 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4903 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4904 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4905 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4906 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4907 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4908 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4909 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4910 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4911 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4912 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4913 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4914 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4915 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4916 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4917 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4918 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4919 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4920 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4921 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4922 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4923 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4924 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4925 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4926 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4927 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4928 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4929 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4930 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4931 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4932 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4933 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4934 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4935 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4936 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4937 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4938 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4939 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4940 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4941 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4942 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4943 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4944 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4945 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4946 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4947 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4948 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4949 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4950 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4951 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4952 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4953 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4954 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4955 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4956 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4957 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4958 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4959 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4960 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4961 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4962 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4963 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4964 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4965 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4966 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4967 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4968 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4969 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4970 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4971 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4972 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4973 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4974 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4975 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4976 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4977 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4978 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4979 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4980 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4981 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4982 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4983 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4984 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4985 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4986 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4987 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4988 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4989 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4990 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4991 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4992 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4993 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4994 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4995 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4996 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4997 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4998 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		4999 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5000 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5001 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5002 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5003 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5004 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5005 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5006 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5007 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5008 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5009 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5010 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5011 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5012 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5013 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5014 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5015 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5016 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5017 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5018 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5019 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5020 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5021 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5022 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5023 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5024 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5025 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5026 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5027 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5028 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5029 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5030 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5031 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5032 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5033 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5034 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5035 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5036 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5037 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5038 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5039 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5040 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5041 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5042 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5043 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5044 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5045 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5046 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5047 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5048 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5049 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5050 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5051 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5052 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5053 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5054 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5055 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5056 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5057 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5058 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5059 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5060 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5061 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5062 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5063 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5064 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5065 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5066 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5067 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5068 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5069 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5070 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5071 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5072 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5073 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5074 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5075 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5076 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5077 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5078 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5079 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5080 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5081 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5082 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5083 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5084 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5085 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5086 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5087 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5088 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5089 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5090 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5091 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5092 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5093 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5094 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5095 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5096 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5097 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5098 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5099 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5100 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5101 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5102 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5103 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5104 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5105 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5106 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5107 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5108 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5109 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5110 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5111 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5112 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5113 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5114 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5115 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5116 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5117 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5118 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5119 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5120 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5121 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5122 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5123 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5124 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5125 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5126 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5127 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5128 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5129 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5130 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5131 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5132 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5133 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5134 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5135 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5136 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5137 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5138 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5139 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5140 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5141 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5142 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5143 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5144 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5145 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5146 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5147 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5148 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5149 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5150 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5151 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5152 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5153 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5154 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5155 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5156 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5157 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5158 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5159 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5160 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5161 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5162 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5163 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5164 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5165 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5166 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5167 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5168 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5169 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5170 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5171 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5172 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5173 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5174 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5175 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5176 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5177 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5178 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5179 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5180 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5181 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5182 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5183 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5184 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5185 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5186 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5187 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5188 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5189 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5190 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5191 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5192 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5193 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5194 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5195 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5196 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5197 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5198 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5199 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5200 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5201 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5202 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5203 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5204 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5205 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5206 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5207 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5208 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5209 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5210 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5211 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5212 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5213 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5214 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5215 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5216 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5217 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5218 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5219 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5220 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5221 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5222 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5223 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5224 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5225 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5226 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5227 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5228 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5229 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5230 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5231 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5232 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5233 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5234 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5235 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5236 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5237 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5238 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5239 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5240 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5241 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5242 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5243 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5244 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5245 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5246 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5247 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5248 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5249 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5250 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5251 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5252 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5253 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5254 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5255 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5256 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5257 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5258 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5259 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5260 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5261 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5262 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5263 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5264 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5265 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5266 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5267 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5268 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5269 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5270 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5271 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5272 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5273 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5274 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5275 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5276 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5277 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5278 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5279 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5280 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5281 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5282 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5283 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5284 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5285 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5286 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5287 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5288 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5289 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5290 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5291 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5292 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5293 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5294 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5295 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5296 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5297 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5298 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5299 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5300 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5301 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5302 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5303 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5304 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5305 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5306 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5307 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5308 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5309 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5310 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5311 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5312 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5313 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5314 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5315 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5316 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5317 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5318 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5319 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5320 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5321 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5322 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5323 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5324 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5325 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5326 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5327 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5328 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5329 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5330 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5331 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5332 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5333 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5334 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5335 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5336 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5337 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5338 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5339 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5340 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5341 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5342 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5343 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5344 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5345 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5346 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5347 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5348 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5349 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5350 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5351 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5352 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5353 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5354 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5355 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5356 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5357 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5358 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5359 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5360 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5361 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5362 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5363 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5364 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5365 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5366 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5367 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5368 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5369 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5370 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5371 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5372 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5373 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5374 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5375 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5376 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5377 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5378 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5379 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5380 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5381 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5382 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5383 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5384 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5385 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5386 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5387 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5388 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5389 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5390 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5391 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5392 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5393 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5394 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5395 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5396 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5397 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5398 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5399 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5400 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5401 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5402 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5403 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5404 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5405 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5406 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5407 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5408 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5409 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5410 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5411 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5412 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5413 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5414 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5415 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5416 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5417 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5418 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5419 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5420 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5421 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5422 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5423 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5424 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5425 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5426 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5427 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5428 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5429 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5430 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5431 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5432 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5433 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5434 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5435 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5436 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5437 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5438 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5439 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5440 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5441 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5442 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5443 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5444 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5445 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5446 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5447 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5448 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5449 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5450 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5451 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5452 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5453 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5454 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5455 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5456 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5457 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5458 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5459 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5460 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5461 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5462 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5463 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5464 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5465 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5466 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5467 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5468 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5469 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5470 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5471 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5472 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5473 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5474 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5475 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5476 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5477 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5478 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5479 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5480 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5481 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5482 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5483 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5484 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5485 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5486 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5487 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5488 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5489 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5490 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5491 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5492 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5493 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5494 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5495 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5496 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5497 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5498 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5499 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5500 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5501 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5502 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5503 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5504 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5505 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5506 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5507 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5508 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5509 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5510 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5511 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5512 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5513 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5514 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5515 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5516 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5517 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5518 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5519 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5520 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5521 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5522 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5523 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5524 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5525 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5526 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5527 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5528 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5529 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5530 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5531 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5532 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5533 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5534 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5535 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5536 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5537 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5538 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5539 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5540 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5541 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5542 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5543 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5544 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5545 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5546 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5547 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5548 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5549 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5550 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5551 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5552 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5553 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5554 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5555 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5556 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5557 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5558 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5559 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5560 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5561 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5562 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5563 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5564 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5565 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5566 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5567 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5568 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5569 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5570 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5571 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5572 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5573 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5574 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5575 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5576 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5577 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5578 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5579 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5580 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5581 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5582 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5583 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5584 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5585 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5586 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5587 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5588 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5589 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5590 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5591 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5592 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5593 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5594 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5595 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5596 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5597 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5598 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5599 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5600 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5601 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5602 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5603 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5604 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5605 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5606 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5607 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5608 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5609 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5610 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5611 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5612 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5613 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5614 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5615 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5616 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5617 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5618 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5619 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5620 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5621 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5622 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5623 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5624 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5625 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5626 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5627 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5628 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5629 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5630 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5631 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5632 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5633 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5634 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5635 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5636 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5637 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5638 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5639 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5640 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5641 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5642 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5643 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5644 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5645 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5646 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5647 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5648 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5649 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5650 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5651 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5652 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5653 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5654 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5655 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5656 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5657 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5658 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5659 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5660 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5661 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5662 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5663 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5664 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5665 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5666 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5667 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5668 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5669 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5670 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5671 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5672 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5673 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5674 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5675 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5676 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5677 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5678 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5679 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5680 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5681 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5682 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5683 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5684 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5685 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5686 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5687 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5688 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5689 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5690 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5691 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5692 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5693 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5694 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5695 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5696 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5697 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5698 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5699 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5700 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5701 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5702 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5703 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5704 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5705 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5706 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5707 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5708 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5709 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5710 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5711 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5712 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5713 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5714 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5715 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5716 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5717 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5718 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5719 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5720 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5721 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5722 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5723 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5724 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5725 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5726 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5727 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5728 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5729 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5730 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5731 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5732 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5733 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5734 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5735 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5736 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5737 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5738 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5739 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5740 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5741 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5742 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5743 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5744 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5745 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5746 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5747 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5748 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5749 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5750 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5751 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5752 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5753 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5754 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5755 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5756 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5757 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5758 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5759 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5760 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5761 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5762 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5763 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5764 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5765 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5766 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5767 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5768 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5769 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5770 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5771 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5772 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5773 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5774 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5775 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5776 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5777 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5778 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5779 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5780 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5781 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5782 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5783 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5784 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5785 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5786 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5787 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5788 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5789 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5790 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5791 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5792 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5793 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5794 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5795 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5796 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5797 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5798 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5799 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5800 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5801 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5802 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5803 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5804 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5805 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5806 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5807 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5808 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5809 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5810 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5811 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5812 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5813 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5814 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5815 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5816 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5817 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5818 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5819 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5820 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5821 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5822 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5823 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5824 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5825 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5826 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5827 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5828 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5829 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5830 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5831 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5832 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5833 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5834 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5835 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5836 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5837 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5838 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5839 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5840 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5841 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5842 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5843 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5844 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5845 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5846 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5847 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5848 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5849 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5850 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5851 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5852 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5853 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5854 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5855 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5856 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5857 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5858 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5859 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5860 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5861 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5862 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5863 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5864 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5865 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5866 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5867 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5868 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5869 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5870 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5871 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5872 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5873 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5874 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5875 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5876 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5877 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5878 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5879 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5880 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5881 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5882 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5883 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5884 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5885 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5886 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5887 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5888 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5889 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5890 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5891 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5892 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5893 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5894 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5895 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5896 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5897 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5898 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5899 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5900 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5901 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5902 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5903 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5904 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5905 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5906 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5907 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5908 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5909 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5910 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5911 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5912 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5913 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5914 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5915 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5916 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5917 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5918 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5919 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5920 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5921 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5922 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5923 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5924 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5925 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5926 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5927 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5928 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5929 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5930 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5931 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5932 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5933 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5934 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5935 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5936 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5937 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5938 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5939 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5940 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5941 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5942 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5943 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5944 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5945 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5946 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5947 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5948 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5949 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5950 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5951 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5952 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5953 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5954 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5955 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5956 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5957 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5958 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5959 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5960 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5961 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5962 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5963 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5964 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5965 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5966 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5967 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5968 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5969 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5970 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5971 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5972 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5973 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5974 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5975 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5976 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5977 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5978 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5979 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5980 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5981 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5982 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5983 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5984 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5985 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5986 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5987 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5988 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5989 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5990 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5991 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5992 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5993 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5994 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5995 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5996 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5997 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5998 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		5999 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6000 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6001 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6002 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6003 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6004 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6005 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6006 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6007 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6008 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6009 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6010 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6011 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6012 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6013 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6014 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6015 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6016 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6017 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6018 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6019 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6020 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6021 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6022 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6023 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6024 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6025 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6026 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6027 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6028 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6029 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6030 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6031 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6032 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6033 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6034 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6035 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6036 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6037 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6038 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6039 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6040 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6041 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6042 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6043 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6044 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6045 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6046 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6047 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6048 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6049 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6050 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6051 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6052 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6053 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6054 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6055 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6056 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6057 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6058 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6059 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6060 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6061 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6062 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6063 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6064 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6065 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6066 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6067 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6068 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6069 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6070 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6071 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6072 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6073 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6074 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6075 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6076 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6077 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6078 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6079 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6080 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6081 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6082 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6083 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6084 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6085 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6086 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6087 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6088 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6089 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6090 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6091 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6092 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6093 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6094 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6095 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6096 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6097 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6098 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6099 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6100 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6101 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6102 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6103 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6104 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6105 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6106 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6107 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6108 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6109 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6110 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6111 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6112 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6113 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6114 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6115 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6116 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6117 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6118 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6119 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6120 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6121 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6122 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6123 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6124 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6125 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6126 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6127 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6128 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6129 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6130 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6131 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6132 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6133 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6134 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6135 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6136 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6137 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6138 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6139 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6140 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6141 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6142 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6143 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6144 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6145 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6146 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6147 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6148 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6149 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6150 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6151 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6152 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6153 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6154 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6155 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6156 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6157 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6158 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6159 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6160 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6161 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6162 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6163 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6164 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6165 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6166 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6167 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6168 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6169 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6170 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6171 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6172 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6173 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6174 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6175 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6176 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6177 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6178 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6179 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6180 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6181 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6182 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6183 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6184 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6185 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6186 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6187 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6188 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6189 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6190 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6191 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6192 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6193 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6194 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6195 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6196 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6197 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6198 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6199 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6200 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6201 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6202 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6203 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6204 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6205 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6206 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6207 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6208 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6209 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6210 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6211 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6212 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6213 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6214 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6215 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6216 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6217 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6218 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6219 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6220 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6221 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6222 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		6223 =>	"00000000000000000000000101100000", -- z: 0 rot: 0 ptr: 352
		others => "00000000000000000000000000000000"
	);

begin

	process( clk_i, mem, addr_i ) begin
		if rising_edge( clk_i ) then
--			if we_i = '1' then
--				mem( to_integer( unsigned( addr_i ) ) ) <= data_o;
--			else
				data_o <= mem( to_integer( unsigned( addr_i ) ) );
--			end if;
		end if; 
	end process;

end architecture arch;