
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);
	
	port
	(
		clk_i    : in  	std_logic;
		addr_i	: in  	std_logic_vector( ADDR_WIDTH-1 downto 0 );
		data_o	: out	std_logic_vector( DATA_WIDTH-1 downto 0 )
	);
end entity ram;

architecture arch of ram is

	type	ram_t is array ( 0 to 2**ADDR_WIDTH-1 ) of std_logic_vector( DATA_WIDTH-1 downto 0 );
	
-- GENERATED BY BC_MEM_PACKER
-- DATE: Sun May 24 17:03:19 2015

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


		0 =>	"10000000000000000000000000000000", -- R: 128 G: 0 B: 0
		1 =>	"01100000011000001000000000000000", -- R: 96 G: 96 B: 128
		2 =>	"10100000010000000000000000000000", -- R: 160 G: 64 B: 0
		3 =>	"00000000000000000000000000000000", -- R: 0 G: 0 B: 0
		4 =>	"10100000101000001010010000000000", -- R: 160 G: 160 B: 164
		5 =>	"00000000011000000000000000000000", -- R: 0 G: 96 B: 0
		6 =>	"00000000010000000000000000000000", -- R: 0 G: 64 B: 0
		7 =>	"10000000111000000000000000000000", -- R: 128 G: 224 B: 0
		8 =>	"11111111111111111111111100000000", -- R: 255 G: 255 B: 255
		9 =>	"01000000010000001100000000000000", -- R: 64 G: 64 B: 192
		10 =>	"10100110110010101111000000000000", -- R: 166 G: 202 B: 240
		11 =>	"00000000010000000100000000000000", -- R: 0 G: 64 B: 64
		12 =>	"01100000000000001000000000000000", -- R: 96 G: 0 B: 128
		13 =>	"11000000010000000100000000000000", -- R: 192 G: 64 B: 64
		14 =>	"11100000111000001000000000000000", -- R: 224 G: 224 B: 128
		15 =>	"11100000101000000100000000000000", -- R: 224 G: 160 B: 64
		16 =>	"01100000011000000000000000000000", -- R: 96 G: 96 B: 0
		17 =>	"00000000000000000000000000000000", -- Unused
		18 =>	"00000000000000000000000000000000", -- Unused
		19 =>	"00000000000000000000000000000000", -- Unused
		20 =>	"00000000000000000000000000000000", -- Unused
		21 =>	"00000000000000000000000000000000", -- Unused
		22 =>	"00000000000000000000000000000000", -- Unused
		23 =>	"00000000000000000000000000000000", -- Unused
		24 =>	"00000000000000000000000000000000", -- Unused
		25 =>	"00000000000000000000000000000000", -- Unused
		26 =>	"00000000000000000000000000000000", -- Unused
		27 =>	"00000000000000000000000000000000", -- Unused
		28 =>	"00000000000000000000000000000000", -- Unused
		29 =>	"00000000000000000000000000000000", -- Unused
		30 =>	"00000000000000000000000000000000", -- Unused
		31 =>	"00000000000000000000000000000000", -- Unused
		32 =>	"00000000000000000000000000000000", -- Unused
		33 =>	"00000000000000000000000000000000", -- Unused
		34 =>	"00000000000000000000000000000000", -- Unused
		35 =>	"00000000000000000000000000000000", -- Unused
		36 =>	"00000000000000000000000000000000", -- Unused
		37 =>	"00000000000000000000000000000000", -- Unused
		38 =>	"00000000000000000000000000000000", -- Unused
		39 =>	"00000000000000000000000000000000", -- Unused
		40 =>	"00000000000000000000000000000000", -- Unused
		41 =>	"00000000000000000000000000000000", -- Unused
		42 =>	"00000000000000000000000000000000", -- Unused
		43 =>	"00000000000000000000000000000000", -- Unused
		44 =>	"00000000000000000000000000000000", -- Unused
		45 =>	"00000000000000000000000000000000", -- Unused
		46 =>	"00000000000000000000000000000000", -- Unused
		47 =>	"00000000000000000000000000000000", -- Unused
		48 =>	"00000000000000000000000000000000", -- Unused
		49 =>	"00000000000000000000000000000000", -- Unused
		50 =>	"00000000000000000000000000000000", -- Unused
		51 =>	"00000000000000000000000000000000", -- Unused
		52 =>	"00000000000000000000000000000000", -- Unused
		53 =>	"00000000000000000000000000000000", -- Unused
		54 =>	"00000000000000000000000000000000", -- Unused
		55 =>	"00000000000000000000000000000000", -- Unused
		56 =>	"00000000000000000000000000000000", -- Unused
		57 =>	"00000000000000000000000000000000", -- Unused
		58 =>	"00000000000000000000000000000000", -- Unused
		59 =>	"00000000000000000000000000000000", -- Unused
		60 =>	"00000000000000000000000000000000", -- Unused
		61 =>	"00000000000000000000000000000000", -- Unused
		62 =>	"00000000000000000000000000000000", -- Unused
		63 =>	"00000000000000000000000000000000", -- Unused
		64 =>	"00000000000000000000000000000000", -- Unused
		65 =>	"00000000000000000000000000000000", -- Unused
		66 =>	"00000000000000000000000000000000", -- Unused
		67 =>	"00000000000000000000000000000000", -- Unused
		68 =>	"00000000000000000000000000000000", -- Unused
		69 =>	"00000000000000000000000000000000", -- Unused
		70 =>	"00000000000000000000000000000000", -- Unused
		71 =>	"00000000000000000000000000000000", -- Unused
		72 =>	"00000000000000000000000000000000", -- Unused
		73 =>	"00000000000000000000000000000000", -- Unused
		74 =>	"00000000000000000000000000000000", -- Unused
		75 =>	"00000000000000000000000000000000", -- Unused
		76 =>	"00000000000000000000000000000000", -- Unused
		77 =>	"00000000000000000000000000000000", -- Unused
		78 =>	"00000000000000000000000000000000", -- Unused
		79 =>	"00000000000000000000000000000000", -- Unused
		80 =>	"00000000000000000000000000000000", -- Unused
		81 =>	"00000000000000000000000000000000", -- Unused
		82 =>	"00000000000000000000000000000000", -- Unused
		83 =>	"00000000000000000000000000000000", -- Unused
		84 =>	"00000000000000000000000000000000", -- Unused
		85 =>	"00000000000000000000000000000000", -- Unused
		86 =>	"00000000000000000000000000000000", -- Unused
		87 =>	"00000000000000000000000000000000", -- Unused
		88 =>	"00000000000000000000000000000000", -- Unused
		89 =>	"00000000000000000000000000000000", -- Unused
		90 =>	"00000000000000000000000000000000", -- Unused
		91 =>	"00000000000000000000000000000000", -- Unused
		92 =>	"00000000000000000000000000000000", -- Unused
		93 =>	"00000000000000000000000000000000", -- Unused
		94 =>	"00000000000000000000000000000000", -- Unused
		95 =>	"00000000000000000000000000000000", -- Unused
		96 =>	"00000000000000000000000000000000", -- Unused
		97 =>	"00000000000000000000000000000000", -- Unused
		98 =>	"00000000000000000000000000000000", -- Unused
		99 =>	"00000000000000000000000000000000", -- Unused
		100 =>	"00000000000000000000000000000000", -- Unused
		101 =>	"00000000000000000000000000000000", -- Unused
		102 =>	"00000000000000000000000000000000", -- Unused
		103 =>	"00000000000000000000000000000000", -- Unused
		104 =>	"00000000000000000000000000000000", -- Unused
		105 =>	"00000000000000000000000000000000", -- Unused
		106 =>	"00000000000000000000000000000000", -- Unused
		107 =>	"00000000000000000000000000000000", -- Unused
		108 =>	"00000000000000000000000000000000", -- Unused
		109 =>	"00000000000000000000000000000000", -- Unused
		110 =>	"00000000000000000000000000000000", -- Unused
		111 =>	"00000000000000000000000000000000", -- Unused
		112 =>	"00000000000000000000000000000000", -- Unused
		113 =>	"00000000000000000000000000000000", -- Unused
		114 =>	"00000000000000000000000000000000", -- Unused
		115 =>	"00000000000000000000000000000000", -- Unused
		116 =>	"00000000000000000000000000000000", -- Unused
		117 =>	"00000000000000000000000000000000", -- Unused
		118 =>	"00000000000000000000000000000000", -- Unused
		119 =>	"00000000000000000000000000000000", -- Unused
		120 =>	"00000000000000000000000000000000", -- Unused
		121 =>	"00000000000000000000000000000000", -- Unused
		122 =>	"00000000000000000000000000000000", -- Unused
		123 =>	"00000000000000000000000000000000", -- Unused
		124 =>	"00000000000000000000000000000000", -- Unused
		125 =>	"00000000000000000000000000000000", -- Unused
		126 =>	"00000000000000000000000000000000", -- Unused
		127 =>	"00000000000000000000000000000000", -- Unused
		128 =>	"00000000000000000000000000000000", -- Unused
		129 =>	"00000000000000000000000000000000", -- Unused
		130 =>	"00000000000000000000000000000000", -- Unused
		131 =>	"00000000000000000000000000000000", -- Unused
		132 =>	"00000000000000000000000000000000", -- Unused
		133 =>	"00000000000000000000000000000000", -- Unused
		134 =>	"00000000000000000000000000000000", -- Unused
		135 =>	"00000000000000000000000000000000", -- Unused
		136 =>	"00000000000000000000000000000000", -- Unused
		137 =>	"00000000000000000000000000000000", -- Unused
		138 =>	"00000000000000000000000000000000", -- Unused
		139 =>	"00000000000000000000000000000000", -- Unused
		140 =>	"00000000000000000000000000000000", -- Unused
		141 =>	"00000000000000000000000000000000", -- Unused
		142 =>	"00000000000000000000000000000000", -- Unused
		143 =>	"00000000000000000000000000000000", -- Unused
		144 =>	"00000000000000000000000000000000", -- Unused
		145 =>	"00000000000000000000000000000000", -- Unused
		146 =>	"00000000000000000000000000000000", -- Unused
		147 =>	"00000000000000000000000000000000", -- Unused
		148 =>	"00000000000000000000000000000000", -- Unused
		149 =>	"00000000000000000000000000000000", -- Unused
		150 =>	"00000000000000000000000000000000", -- Unused
		151 =>	"00000000000000000000000000000000", -- Unused
		152 =>	"00000000000000000000000000000000", -- Unused
		153 =>	"00000000000000000000000000000000", -- Unused
		154 =>	"00000000000000000000000000000000", -- Unused
		155 =>	"00000000000000000000000000000000", -- Unused
		156 =>	"00000000000000000000000000000000", -- Unused
		157 =>	"00000000000000000000000000000000", -- Unused
		158 =>	"00000000000000000000000000000000", -- Unused
		159 =>	"00000000000000000000000000000000", -- Unused
		160 =>	"00000000000000000000000000000000", -- Unused
		161 =>	"00000000000000000000000000000000", -- Unused
		162 =>	"00000000000000000000000000000000", -- Unused
		163 =>	"00000000000000000000000000000000", -- Unused
		164 =>	"00000000000000000000000000000000", -- Unused
		165 =>	"00000000000000000000000000000000", -- Unused
		166 =>	"00000000000000000000000000000000", -- Unused
		167 =>	"00000000000000000000000000000000", -- Unused
		168 =>	"00000000000000000000000000000000", -- Unused
		169 =>	"00000000000000000000000000000000", -- Unused
		170 =>	"00000000000000000000000000000000", -- Unused
		171 =>	"00000000000000000000000000000000", -- Unused
		172 =>	"00000000000000000000000000000000", -- Unused
		173 =>	"00000000000000000000000000000000", -- Unused
		174 =>	"00000000000000000000000000000000", -- Unused
		175 =>	"00000000000000000000000000000000", -- Unused
		176 =>	"00000000000000000000000000000000", -- Unused
		177 =>	"00000000000000000000000000000000", -- Unused
		178 =>	"00000000000000000000000000000000", -- Unused
		179 =>	"00000000000000000000000000000000", -- Unused
		180 =>	"00000000000000000000000000000000", -- Unused
		181 =>	"00000000000000000000000000000000", -- Unused
		182 =>	"00000000000000000000000000000000", -- Unused
		183 =>	"00000000000000000000000000000000", -- Unused
		184 =>	"00000000000000000000000000000000", -- Unused
		185 =>	"00000000000000000000000000000000", -- Unused
		186 =>	"00000000000000000000000000000000", -- Unused
		187 =>	"00000000000000000000000000000000", -- Unused
		188 =>	"00000000000000000000000000000000", -- Unused
		189 =>	"00000000000000000000000000000000", -- Unused
		190 =>	"00000000000000000000000000000000", -- Unused
		191 =>	"00000000000000000000000000000000", -- Unused
		192 =>	"00000000000000000000000000000000", -- Unused
		193 =>	"00000000000000000000000000000000", -- Unused
		194 =>	"00000000000000000000000000000000", -- Unused
		195 =>	"00000000000000000000000000000000", -- Unused
		196 =>	"00000000000000000000000000000000", -- Unused
		197 =>	"00000000000000000000000000000000", -- Unused
		198 =>	"00000000000000000000000000000000", -- Unused
		199 =>	"00000000000000000000000000000000", -- Unused
		200 =>	"00000000000000000000000000000000", -- Unused
		201 =>	"00000000000000000000000000000000", -- Unused
		202 =>	"00000000000000000000000000000000", -- Unused
		203 =>	"00000000000000000000000000000000", -- Unused
		204 =>	"00000000000000000000000000000000", -- Unused
		205 =>	"00000000000000000000000000000000", -- Unused
		206 =>	"00000000000000000000000000000000", -- Unused
		207 =>	"00000000000000000000000000000000", -- Unused
		208 =>	"00000000000000000000000000000000", -- Unused
		209 =>	"00000000000000000000000000000000", -- Unused
		210 =>	"00000000000000000000000000000000", -- Unused
		211 =>	"00000000000000000000000000000000", -- Unused
		212 =>	"00000000000000000000000000000000", -- Unused
		213 =>	"00000000000000000000000000000000", -- Unused
		214 =>	"00000000000000000000000000000000", -- Unused
		215 =>	"00000000000000000000000000000000", -- Unused
		216 =>	"00000000000000000000000000000000", -- Unused
		217 =>	"00000000000000000000000000000000", -- Unused
		218 =>	"00000000000000000000000000000000", -- Unused
		219 =>	"00000000000000000000000000000000", -- Unused
		220 =>	"00000000000000000000000000000000", -- Unused
		221 =>	"00000000000000000000000000000000", -- Unused
		222 =>	"00000000000000000000000000000000", -- Unused
		223 =>	"00000000000000000000000000000000", -- Unused
		224 =>	"00000000000000000000000000000000", -- Unused
		225 =>	"00000000000000000000000000000000", -- Unused
		226 =>	"00000000000000000000000000000000", -- Unused
		227 =>	"00000000000000000000000000000000", -- Unused
		228 =>	"00000000000000000000000000000000", -- Unused
		229 =>	"00000000000000000000000000000000", -- Unused
		230 =>	"00000000000000000000000000000000", -- Unused
		231 =>	"00000000000000000000000000000000", -- Unused
		232 =>	"00000000000000000000000000000000", -- Unused
		233 =>	"00000000000000000000000000000000", -- Unused
		234 =>	"00000000000000000000000000000000", -- Unused
		235 =>	"00000000000000000000000000000000", -- Unused
		236 =>	"00000000000000000000000000000000", -- Unused
		237 =>	"00000000000000000000000000000000", -- Unused
		238 =>	"00000000000000000000000000000000", -- Unused
		239 =>	"00000000000000000000000000000000", -- Unused
		240 =>	"00000000000000000000000000000000", -- Unused
		241 =>	"00000000000000000000000000000000", -- Unused
		242 =>	"00000000000000000000000000000000", -- Unused
		243 =>	"00000000000000000000000000000000", -- Unused
		244 =>	"00000000000000000000000000000000", -- Unused
		245 =>	"00000000000000000000000000000000", -- Unused
		246 =>	"00000000000000000000000000000000", -- Unused
		247 =>	"00000000000000000000000000000000", -- Unused
		248 =>	"00000000000000000000000000000000", -- Unused
		249 =>	"00000000000000000000000000000000", -- Unused
		250 =>	"00000000000000000000000000000000", -- Unused
		251 =>	"00000000000000000000000000000000", -- Unused
		252 =>	"00000000000000000000000000000000", -- Unused
		253 =>	"00000000000000000000000000000000", -- Unused
		254 =>	"00000000000000000000000000000000", -- Unused
		255 =>	"00000000000000000000000000000000", -- Unused


--			***** 8x8 IMAGES *****


		256 =>	"00000000000000000000000000000000", -- IMG_8x8_BRICK
		257 =>	"00000001000000000000000000000000",
		258 =>	"00000010000000100000001000000010",
		259 =>	"00000001000000000000001000000010",
		260 =>	"00000010000000100000001000000010",
		261 =>	"00000001000000000000001000000010",
		262 =>	"00000001000000010000000100000001",
		263 =>	"00000001000000010000000100000001",
		264 =>	"00000001000000000000000000000000",
		265 =>	"00000000000000000000000000000000",
		266 =>	"00000001000000000000001000000010",
		267 =>	"00000010000000100000001000000010",
		268 =>	"00000001000000000000001000000010",
		269 =>	"00000010000000100000001000000010",
		270 =>	"00000001000000010000000100000001",
		271 =>	"00000001000000010000000100000001",
		272 =>	"00000011000000110000001100000011", -- IMG_8x8_BULLET
		273 =>	"00000011000000110000001100000011",
		274 =>	"00000011000000110000001100000011",
		275 =>	"00000011000000110000001100000011",
		276 =>	"00000011000000110000001100000100",
		277 =>	"00000011000000110000001100000011",
		278 =>	"00000011000000110000010000000100",
		279 =>	"00000100000000110000001100000011",
		280 =>	"00000011000000110000010000000100",
		281 =>	"00000100000000110000001100000011",
		282 =>	"00000011000000110000010000000100",
		283 =>	"00000100000000110000001100000011",
		284 =>	"00000011000000110000001100000011",
		285 =>	"00000011000000110000001100000011",
		286 =>	"00000011000000110000001100000011",
		287 =>	"00000011000000110000001100000011",
		288 =>	"00000011000001010000010100000101", -- IMG_8x8_GRASS
		289 =>	"00000110000001010000011100000011",
		290 =>	"00000101000001010000011000000111",
		291 =>	"00000101000001110000010100000111",
		292 =>	"00000101000001010000010100000101",
		293 =>	"00000101000001110000011100000111",
		294 =>	"00000110000001010000010100000111",
		295 =>	"00000111000001100000010100000111",
		296 =>	"00000101000001010000011100000110",
		297 =>	"00000111000001110000011100000110",
		298 =>	"00000101000001100000010100000111",
		299 =>	"00000111000001110000011100000111",
		300 =>	"00000111000001110000011100000111",
		301 =>	"00000111000001100000011100000111",
		302 =>	"00000011000001110000011100000110",
		303 =>	"00000111000001110000011100000011",
		304 =>	"00000001000001000000010000001000", -- IMG_8x8_ICE
		305 =>	"00000001000001000000010000001000",
		306 =>	"00000100000001000000010000000100",
		307 =>	"00000100000001000000100000000001",
		308 =>	"00000100000001000000010000000100",
		309 =>	"00000100000010000000000100000100",
		310 =>	"00001000000001000000010000000100",
		311 =>	"00001000000000010000010000000100",
		312 =>	"00000001000001000000010000001000",
		313 =>	"00000001000001000000010000001000",
		314 =>	"00000100000001000000100000000001",
		315 =>	"00000100000001000000100000000001",
		316 =>	"00000100000010000000000100000100",
		317 =>	"00000100000010000000000100000100",
		318 =>	"00001000000000010000010000000100",
		319 =>	"00001000000000010000010000000100",
		320 =>	"00000100000001000000010000000100", -- IMG_8x8_IRON
		321 =>	"00000100000001000000010000000100",
		322 =>	"00000100000001000000010000000100",
		323 =>	"00000100000001000000010000000001",
		324 =>	"00000100000001000000100000001000",
		325 =>	"00001000000010000000000100000001",
		326 =>	"00000100000001000000100000001000",
		327 =>	"00001000000010000000000100000001",
		328 =>	"00000100000001000000100000001000",
		329 =>	"00001000000010000000000100000001",
		330 =>	"00000100000001000000100000001000",
		331 =>	"00001000000010000000000100000001",
		332 =>	"00000100000001000000000100000001",
		333 =>	"00000001000000010000000100000001",
		334 =>	"00000100000000010000000100000001",
		335 =>	"00000001000000010000000100000001",
		336 =>	"00000001000000010000000100000010", -- IMG_8x8_LIVES_REMAINING_ICON
		337 =>	"00000010000000100000000100000001",
		338 =>	"00000001000000100000000100000001",
		339 =>	"00000010000000010000000100000010",
		340 =>	"00000001000000100000000100000010",
		341 =>	"00000010000000100000000100000010",
		342 =>	"00000001000000100000001000000010",
		343 =>	"00000001000000100000001000000010",
		344 =>	"00000001000000100000001000000001",
		345 =>	"00000001000000010000001000000010",
		346 =>	"00000001000000100000001000000010",
		347 =>	"00000001000000100000001000000010",
		348 =>	"00000001000000100000000100000010",
		349 =>	"00000010000000100000000100000010",
		350 =>	"00000001000000100000000100000001",
		351 =>	"00000010000000010000000100000010",
		352 =>	"00000001000000010000000100000001", -- IMG_8x8_TANKS_REMAINING_ICON
		353 =>	"00000001000000010000000100000001",
		354 =>	"00000001000000110000000100000001",
		355 =>	"00000011000000010000000100000011",
		356 =>	"00000001000000110000000100000011",
		357 =>	"00000011000000110000000100000011",
		358 =>	"00000001000000110000001100000011",
		359 =>	"00000000000000110000001100000011",
		360 =>	"00000001000000110000001100000011",
		361 =>	"00000000000000110000001100000011",
		362 =>	"00000001000000110000000100000011",
		363 =>	"00000011000000110000000100000011",
		364 =>	"00000001000000110000000100000001",
		365 =>	"00000011000000010000000100000011",
		366 =>	"00000001000000010000000100000011",
		367 =>	"00000011000000110000000100000001",
		368 =>	"00001001000010010000100100001001", -- IMG_8x8_WATER
		369 =>	"00001001000010010000100100001010",
		370 =>	"00001001000010100000100100001001",
		371 =>	"00001001000010010000100100001001",
		372 =>	"00001001000010010000101000001001",
		373 =>	"00001001000010010000100100001001",
		374 =>	"00001001000010010000100100001010",
		375 =>	"00001001000010010000101000001001",
		376 =>	"00001001000010010000100100001001",
		377 =>	"00001001000010010000100100001010",
		378 =>	"00001001000010010000100100001010",
		379 =>	"00001001000010010000100100001001",
		380 =>	"00001001000010010000101000001001",
		381 =>	"00001010000010010000100100001001",
		382 =>	"00001010000010010000100100001001",
		383 =>	"00001001000010010000100100001001",


--			***** 16x16 IMAGES *****


		384 =>	"00000011000000110000001100000011", -- IMG_16x16_BASE_ALIVE
		385 =>	"00000011000000110000001100000011",
		386 =>	"00000011000000110000001100000011",
		387 =>	"00000011000000110000001100000011",
		388 =>	"00000001000000010000001100000011",
		389 =>	"00000011000000110000001100000011",
		390 =>	"00000011000000110000001100000011",
		391 =>	"00000011000000110000000100000001",
		392 =>	"00000011000000010000000100000011",
		393 =>	"00000011000000110000000100000001",
		394 =>	"00000001000000110000001100000011",
		395 =>	"00000011000000010000000100000011",
		396 =>	"00000001000000010000000100000001",
		397 =>	"00000011000000110000001100000001",
		398 =>	"00000000000000010000001100000011",
		399 =>	"00000001000000010000000100000001",
		400 =>	"00000011000000010000000100000001",
		401 =>	"00000011000000110000001100000001",
		402 =>	"00000001000000110000001100000011",
		403 =>	"00000001000000010000000100000011",
		404 =>	"00000001000000010000000100000001",
		405 =>	"00000001000000010000001100000001",
		406 =>	"00000001000000110000000100000001",
		407 =>	"00000001000000010000000100000001",
		408 =>	"00000011000000110000000100000000",
		409 =>	"00000001000000010000000100000001",
		410 =>	"00000001000000010000000100000001",
		411 =>	"00000000000000010000001100000011",
		412 =>	"00000011000000010000000100000001",
		413 =>	"00000000000000010000000100000001",
		414 =>	"00000001000000010000000100000000",
		415 =>	"00000001000000010000000100000011",
		416 =>	"00000011000000110000000100000001",
		417 =>	"00000001000000010000000000000001",
		418 =>	"00000001000000000000000100000001",
		419 =>	"00000001000000010000001100000011",
		420 =>	"00000011000000110000000100000001",
		421 =>	"00000001000000010000000100000001",
		422 =>	"00000001000000010000000100000001",
		423 =>	"00000001000000010000001100000011",
		424 =>	"00000011000000110000001100000001",
		425 =>	"00000001000000010000001100000001",
		426 =>	"00000001000000110000000100000001",
		427 =>	"00000001000000110000001100000011",
		428 =>	"00000011000000110000001100000011",
		429 =>	"00000011000000110000001100000001",
		430 =>	"00000001000000110000001100000011",
		431 =>	"00000011000000110000001100000011",
		432 =>	"00000011000000110000001100000011",
		433 =>	"00000011000000110000000100000001",
		434 =>	"00000001000000010000001100000011",
		435 =>	"00000011000000110000001100000011",
		436 =>	"00000011000000110000001100000011",
		437 =>	"00000001000000010000000100000001",
		438 =>	"00000001000000010000000100000001",
		439 =>	"00000011000000110000001100000011",
		440 =>	"00000011000000110000001100000011",
		441 =>	"00000001000000010000001100000001",
		442 =>	"00000001000000110000000100000001",
		443 =>	"00000011000000110000001100000011",
		444 =>	"00000011000000110000001100000011",
		445 =>	"00000011000000110000001100000011",
		446 =>	"00000011000000110000001100000011",
		447 =>	"00000011000000110000001100000011",
		448 =>	"00000011000000110000001100000011", -- IMG_16x16_BASE_DEAD
		449 =>	"00000011000000110000001100000011",
		450 =>	"00000011000000110000001100000011",
		451 =>	"00000011000000110000001100000011",
		452 =>	"00000011000000110000001100000011",
		453 =>	"00000011000000100000001100000011",
		454 =>	"00000011000000110000001100000011",
		455 =>	"00000011000000110000001100000011",
		456 =>	"00000011000000110000001100000011",
		457 =>	"00000010000000100000001100000001",
		458 =>	"00000011000000110000001100000011",
		459 =>	"00000011000000110000001100000011",
		460 =>	"00000011000000110000001100000011",
		461 =>	"00000010000000110000000100000001",
		462 =>	"00000001000000110000001100000011",
		463 =>	"00000011000000110000001100000011",
		464 =>	"00000011000000110000001100000010",
		465 =>	"00000011000000010000000100000001",
		466 =>	"00000001000000010000001100000011",
		467 =>	"00000011000000110000001100000011",
		468 =>	"00000011000000110000001000000010",
		469 =>	"00000011000000010000000100000001",
		470 =>	"00000001000000010000000100000001",
		471 =>	"00000001000000110000001100000011",
		472 =>	"00000011000000110000001000000011",
		473 =>	"00000001000000010000000100000001",
		474 =>	"00000001000000010000000100000001",
		475 =>	"00000001000000010000001100000011",
		476 =>	"00000011000000100000001000000011",
		477 =>	"00000001000000010000000100000001",
		478 =>	"00000001000000010000000100000001",
		479 =>	"00000001000000010000001100000011",
		480 =>	"00000011000000100000001100000011",
		481 =>	"00000001000000010000000100000001",
		482 =>	"00000001000000010000000100000001",
		483 =>	"00000011000000010000000100000011",
		484 =>	"00000011000000100000001100000001",
		485 =>	"00000001000000010000000100000001",
		486 =>	"00000001000000110000001100000001",
		487 =>	"00000011000000010000000100000011",
		488 =>	"00000011000000100000001100000011",
		489 =>	"00000011000000010000000100000001",
		490 =>	"00000011000000110000001100000011",
		491 =>	"00000011000000010000001100000011",
		492 =>	"00000011000000100000001100000011",
		493 =>	"00000011000000110000001100000001",
		494 =>	"00000011000000110000001100000011",
		495 =>	"00000011000000010000001100000011",
		496 =>	"00000011000000100000001100000011",
		497 =>	"00000011000000110000001100000011",
		498 =>	"00000011000000110000001100000011",
		499 =>	"00000011000000110000001100000011",
		500 =>	"00000011000000100000001100000011",
		501 =>	"00000011000000110000001100000011",
		502 =>	"00000011000000110000001100000011",
		503 =>	"00000011000000110000001100000011",
		504 =>	"00000011000000100000001100000011",
		505 =>	"00000011000000110000001100000011",
		506 =>	"00000011000000110000001100000011",
		507 =>	"00000011000000110000001100000011",
		508 =>	"00000011000000110000001100000011",
		509 =>	"00000011000000110000001100000011",
		510 =>	"00000011000000110000001100000011",
		511 =>	"00000011000000110000001100000011",
		512 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_BOMB
		513 =>	"00000011000000110000001100000011",
		514 =>	"00000011000000110000001100000011",
		515 =>	"00000011000000110000001100000011",
		516 =>	"00000011000010000000100000001000",
		517 =>	"00001000000010000000100000001000",
		518 =>	"00001000000010000000100000001000",
		519 =>	"00001000000010000000010000000011",
		520 =>	"00001000000000110000001100000011",
		521 =>	"00000011000000110000001100000011",
		522 =>	"00000011000000110000001100000011",
		523 =>	"00000011000000110000100000001011",
		524 =>	"00001000000000110000101100001011",
		525 =>	"00001011000010000000100000001000",
		526 =>	"00000100000001000000001100001011",
		527 =>	"00001011000010110000100000001011",
		528 =>	"00001000000000110000101100001011",
		529 =>	"00001011000010000000010000001011",
		530 =>	"00000011000000110000010000000011",
		531 =>	"00001011000010110000100000001011",
		532 =>	"00001000000000110000101100001011",
		533 =>	"00001000000001000000010000000100",
		534 =>	"00001011000000110000001100000100",
		535 =>	"00000011000010110000100000001011",
		536 =>	"00001000000000110000101100001000",
		537 =>	"00000100000010110000100000000100",
		538 =>	"00001011000001000000001100000100",
		539 =>	"00000011000010110000100000001011",
		540 =>	"00001000000000110000101100000100",
		541 =>	"00000011000001000000001100000011",
		542 =>	"00000100000000110000001100000100",
		543 =>	"00000011000010110000100000001011",
		544 =>	"00001000000000110000101100001000",
		545 =>	"00000100000010110000100000000100",
		546 =>	"00001011000001000000001100000100",
		547 =>	"00000011000010110000100000001011",
		548 =>	"00001000000000110000101100000100",
		549 =>	"00000011000001000000001100000011",
		550 =>	"00000100000000110000001100000100",
		551 =>	"00000011000010110000100000001011",
		552 =>	"00001000000000110000101100001000",
		553 =>	"00000100000010110000100000000100",
		554 =>	"00001011000001000000001100000011",
		555 =>	"00001011000010110000100000001011",
		556 =>	"00001000000000110000101100001011",
		557 =>	"00000100000010110000001100000011",
		558 =>	"00000100000000110000101100001011",
		559 =>	"00001011000010110000100000001011",
		560 =>	"00001000000000110000101100001011",
		561 =>	"00001011000010000000010000000100",
		562 =>	"00000011000010110000101100001011",
		563 =>	"00001011000010110000100000001011",
		564 =>	"00001000000000110000101100001011",
		565 =>	"00001011000000110000001100000011",
		566 =>	"00001011000010110000101100001011",
		567 =>	"00001011000010110000100000001011",
		568 =>	"00000100000010000000100000001000",
		569 =>	"00001000000010000000100000001000",
		570 =>	"00001000000010000000100000001000",
		571 =>	"00001000000010000000010000001011",
		572 =>	"00000011000010110000101100001011",
		573 =>	"00001011000010110000101100001011",
		574 =>	"00001011000010110000101100001011",
		575 =>	"00001011000010110000101100000011",
		576 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_GUN
		577 =>	"00000011000000110000001100000011",
		578 =>	"00000011000000110000001100000011",
		579 =>	"00000011000000110000001100000011",
		580 =>	"00000011000010000000100000001000",
		581 =>	"00001000000010000000100000001000",
		582 =>	"00001000000010000000100000001000",
		583 =>	"00001000000010000000010000000011",
		584 =>	"00001000000000110000001100000011",
		585 =>	"00000011000000110000001100000011",
		586 =>	"00000011000000110000001100000011",
		587 =>	"00000011000000110000100000001011",
		588 =>	"00001000000000110000101100001011",
		589 =>	"00001011000010110000101100001011",
		590 =>	"00001011000010110000101100001011",
		591 =>	"00001011000010110000100000001011",
		592 =>	"00001000000000110000101100001000",
		593 =>	"00001011000010110000101100001011",
		594 =>	"00001011000010110000101100001011",
		595 =>	"00001011000010110000100000001011",
		596 =>	"00001000000000110000010000001000",
		597 =>	"00001000000010000000100000001000",
		598 =>	"00001000000010000000010000000011",
		599 =>	"00001011000010110000100000001011",
		600 =>	"00001000000000110000100000000100",
		601 =>	"00000100000001000000010000000100",
		602 =>	"00000100000001000000010000000100",
		603 =>	"00000011000010110000100000001011",
		604 =>	"00001000000000110000001100000100",
		605 =>	"00000100000010110000101100001011",
		606 =>	"00001011000010110000101100000100",
		607 =>	"00000011000010110000100000001011",
		608 =>	"00001000000000110000101100000011",
		609 =>	"00000011000001000000010000001011",
		610 =>	"00000100000001000000010000000100",
		611 =>	"00000100000000110000100000001011",
		612 =>	"00001000000000110000101100001011",
		613 =>	"00001011000000110000010000000011",
		614 =>	"00000011000001000000100000001011",
		615 =>	"00000100000000110000100000001011",
		616 =>	"00001000000000110000101100001011",
		617 =>	"00001011000010110000001100000100",
		618 =>	"00000100000001000000100000001011",
		619 =>	"00000100000000110000100000001011",
		620 =>	"00001000000000110000101100001011",
		621 =>	"00001011000010110000101100000011",
		622 =>	"00000011000001000000101100001011",
		623 =>	"00000100000000110000100000001011",
		624 =>	"00001000000000110000101100001011",
		625 =>	"00001011000010110000101100001011",
		626 =>	"00001011000001000000010000000100",
		627 =>	"00000100000000110000100000001011",
		628 =>	"00001000000000110000101100001011",
		629 =>	"00001011000010110000101100001011",
		630 =>	"00001011000000110000001100000011",
		631 =>	"00000011000010110000100000001011",
		632 =>	"00000100000010000000100000001000",
		633 =>	"00001000000010000000100000001000",
		634 =>	"00001000000010000000100000001000",
		635 =>	"00001000000010000000010000001011",
		636 =>	"00000011000010110000101100001011",
		637 =>	"00001011000010110000101100001011",
		638 =>	"00001011000010110000101100001011",
		639 =>	"00001011000010110000101100000011",
		640 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_SHELL
		641 =>	"00000011000000110000001100000011",
		642 =>	"00000011000000110000001100000011",
		643 =>	"00000011000000110000001100000011",
		644 =>	"00000011000010000000100000001000",
		645 =>	"00001000000010000000100000001000",
		646 =>	"00001000000010000000100000001000",
		647 =>	"00001000000010000000010000000011",
		648 =>	"00001000000000110000001100000011",
		649 =>	"00000011000000110000001100000011",
		650 =>	"00000011000000110000001100000011",
		651 =>	"00000011000000110000100000001011",
		652 =>	"00001000000000110000101100001011",
		653 =>	"00001011000010110000101100001011",
		654 =>	"00001011000010110000101100001011",
		655 =>	"00001011000010110000100000001011",
		656 =>	"00001000000000110000101100001011",
		657 =>	"00001011000010110000101100001011",
		658 =>	"00001011000010110000101100001011",
		659 =>	"00001011000010110000100000001011",
		660 =>	"00001000000000110000101100001011",
		661 =>	"00001011000010000000100000001000",
		662 =>	"00000100000001000000001100001011",
		663 =>	"00001011000010110000100000001011",
		664 =>	"00001000000000110000101100001011",
		665 =>	"00001000000010000000010000000100",
		666 =>	"00000100000001000000010000000011",
		667 =>	"00001011000010110000100000001011",
		668 =>	"00001000000000110000101100001011",
		669 =>	"00001000000001000000010000000100",
		670 =>	"00000100000001000000010000000011",
		671 =>	"00001011000010110000100000001011",
		672 =>	"00001000000000110000101100001011",
		673 =>	"00000100000001000000010000000100",
		674 =>	"00000100000001000000010000000011",
		675 =>	"00001011000010110000100000001011",
		676 =>	"00001000000000110000101100000100",
		677 =>	"00000100000001000000010000000100",
		678 =>	"00000100000001000000010000000011",
		679 =>	"00001011000010110000100000001011",
		680 =>	"00001000000000110000101100000011",
		681 =>	"00000011000000110000001100000011",
		682 =>	"00000100000001000000010000000100",
		683 =>	"00000011000010110000100000001011",
		684 =>	"00001000000000110000101100001011",
		685 =>	"00001011000010110000101100001011",
		686 =>	"00000011000000110000001100000011",
		687 =>	"00000011000010110000100000001011",
		688 =>	"00001000000000110000101100001011",
		689 =>	"00001011000010110000101100001011",
		690 =>	"00001011000010110000101100001011",
		691 =>	"00001011000010110000100000001011",
		692 =>	"00001000000000110000101100001011",
		693 =>	"00001011000010110000101100001011",
		694 =>	"00001011000010110000101100001011",
		695 =>	"00001011000010110000100000001011",
		696 =>	"00000100000010000000100000001000",
		697 =>	"00001000000010000000100000001000",
		698 =>	"00001000000010000000100000001000",
		699 =>	"00001000000010000000010000001011",
		700 =>	"00000011000010110000101100001011",
		701 =>	"00001011000010110000101100001011",
		702 =>	"00001011000010110000101100001011",
		703 =>	"00001011000010110000101100000011",
		704 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_SHOVEL
		705 =>	"00000011000000110000001100000011",
		706 =>	"00000011000000110000001100000011",
		707 =>	"00000011000000110000001100000011",
		708 =>	"00000011000010000000100000001000",
		709 =>	"00001000000010000000100000001000",
		710 =>	"00001000000010000000100000001000",
		711 =>	"00001000000010000000010000000011",
		712 =>	"00001000000000110000001100000011",
		713 =>	"00000011000000110000001100000011",
		714 =>	"00000011000000110000001100000011",
		715 =>	"00000011000000110000100000001011",
		716 =>	"00001000000000110000101100001011",
		717 =>	"00001011000010110000101100001011",
		718 =>	"00001011000010110000100000001011",
		719 =>	"00001011000010110000100000001011",
		720 =>	"00001000000000110000101100001011",
		721 =>	"00001011000010110000101100001011",
		722 =>	"00001011000010110000100000000100",
		723 =>	"00001011000010110000100000001011",
		724 =>	"00001000000000110000101100001011",
		725 =>	"00001011000010110000101100001011",
		726 =>	"00001011000010110000010000000100",
		727 =>	"00000100000010110000100000001011",
		728 =>	"00001000000000110000101100001011",
		729 =>	"00001011000010110000101100001011",
		730 =>	"00001011000010000000001100000011",
		731 =>	"00000011000010110000100000001011",
		732 =>	"00001000000000110000101100001011",
		733 =>	"00001011000010000000101100001011",
		734 =>	"00001000000000110000101100001011",
		735 =>	"00001011000010110000100000001011",
		736 =>	"00001000000000110000101100001011",
		737 =>	"00001000000010000000010000001000",
		738 =>	"00000011000010110000101100001011",
		739 =>	"00001011000010110000100000001011",
		740 =>	"00001000000000110000101100001000",
		741 =>	"00001000000001000000101100000100",
		742 =>	"00000011000010110000101100001011",
		743 =>	"00001011000010110000100000001011",
		744 =>	"00001000000000110000101100001000",
		745 =>	"00000100000010110000010000000100",
		746 =>	"00000100000000110000101100001011",
		747 =>	"00001011000010110000100000001011",
		748 =>	"00001000000000110000101100000100",
		749 =>	"00000100000001000000010000000100",
		750 =>	"00000011000010110000101100001011",
		751 =>	"00001011000010110000100000001011",
		752 =>	"00001000000000110000101100000100",
		753 =>	"00000100000001000000010000000011",
		754 =>	"00001011000010110000101100001011",
		755 =>	"00001011000010110000100000001011",
		756 =>	"00001000000000110000101100000011",
		757 =>	"00000011000000110000001100001011",
		758 =>	"00001011000010110000101100001011",
		759 =>	"00001011000010110000100000001011",
		760 =>	"00000100000010000000100000001000",
		761 =>	"00001000000010000000100000001000",
		762 =>	"00001000000010000000100000001000",
		763 =>	"00001000000010000000010000001011",
		764 =>	"00000011000010110000101100001011",
		765 =>	"00001011000010110000101100001011",
		766 =>	"00001011000010110000101100001011",
		767 =>	"00001011000010110000101100000011",
		768 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_STAR
		769 =>	"00000011000000110000001100000011",
		770 =>	"00000011000000110000001100000011",
		771 =>	"00000011000000110000001100000011",
		772 =>	"00000011000010000000100000001000",
		773 =>	"00001000000010000000100000001000",
		774 =>	"00001000000010000000100000001000",
		775 =>	"00001000000010000000010000000011",
		776 =>	"00001000000000110000001100000011",
		777 =>	"00000011000000110000001100000011",
		778 =>	"00000011000000110000001100000011",
		779 =>	"00000011000000110000100000001011",
		780 =>	"00001000000000110000101100001011",
		781 =>	"00001011000010110000101100001000",
		782 =>	"00000011000010110000101100001011",
		783 =>	"00001011000010110000100000001011",
		784 =>	"00001000000000110000101100001011",
		785 =>	"00001011000010110000100000001000",
		786 =>	"00000100000000110000101100001011",
		787 =>	"00001011000010110000100000001011",
		788 =>	"00001000000000110000101100001011",
		789 =>	"00001011000010110000100000001000",
		790 =>	"00000100000000110000101100001011",
		791 =>	"00001011000010110000100000001011",
		792 =>	"00001000000000110000100000001000",
		793 =>	"00001000000010000000100000000100",
		794 =>	"00000100000010000000100000001000",
		795 =>	"00001000000000110000100000001011",
		796 =>	"00001000000000110000101100000100",
		797 =>	"00000100000001000000100000000100",
		798 =>	"00001000000001000000010000000100",
		799 =>	"00000011000000110000100000001011",
		800 =>	"00001000000000110000101100001011",
		801 =>	"00000100000010000000100000001000",
		802 =>	"00001000000001000000010000000011",
		803 =>	"00000011000010110000100000001011",
		804 =>	"00001000000000110000101100001011",
		805 =>	"00001000000010000000010000000100",
		806 =>	"00001000000010000000010000000011",
		807 =>	"00001011000010110000100000001011",
		808 =>	"00001000000000110000101100000100",
		809 =>	"00001000000001000000010000000011",
		810 =>	"00000100000001000000100000000100",
		811 =>	"00000011000010110000100000001011",
		812 =>	"00001000000000110000101100001000",
		813 =>	"00000100000001000000001100000011",
		814 =>	"00000011000001000000010000001000",
		815 =>	"00000011000010110000100000001011",
		816 =>	"00001000000000110000101100000100",
		817 =>	"00000011000000110000001100001011",
		818 =>	"00001011000000110000001100000100",
		819 =>	"00000011000010110000100000001011",
		820 =>	"00001000000000110000101100000011",
		821 =>	"00000011000010110000101100001011",
		822 =>	"00001011000010110000101100000011",
		823 =>	"00000011000010110000100000001011",
		824 =>	"00000100000010000000100000001000",
		825 =>	"00001000000010000000100000001000",
		826 =>	"00001000000010000000100000001000",
		827 =>	"00001000000010000000010000001011",
		828 =>	"00000011000010110000101100001011",
		829 =>	"00001011000010110000101100001011",
		830 =>	"00001011000010110000101100001011",
		831 =>	"00001011000010110000101100000011",
		832 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_TANK
		833 =>	"00000011000000110000001100000011",
		834 =>	"00000011000000110000001100000011",
		835 =>	"00000011000000110000001100000011",
		836 =>	"00000011000010000000100000001000",
		837 =>	"00001000000010000000100000001000",
		838 =>	"00001000000010000000100000001000",
		839 =>	"00001000000010000000010000000011",
		840 =>	"00001000000000110000001100000011",
		841 =>	"00000011000000110000001100000011",
		842 =>	"00000011000000110000001100000011",
		843 =>	"00000011000000110000100000001011",
		844 =>	"00001000000000110000101100001011",
		845 =>	"00001011000010110000101100001011",
		846 =>	"00001011000010110000101100001011",
		847 =>	"00001011000010110000100000001011",
		848 =>	"00001000000000110000101100001000",
		849 =>	"00001011000010110000101100001011",
		850 =>	"00001011000010110000101100001011",
		851 =>	"00001011000010110000100000001011",
		852 =>	"00001000000000110000010000001000",
		853 =>	"00001000000010000000100000001000",
		854 =>	"00001000000010000000010000000011",
		855 =>	"00001011000010110000100000001011",
		856 =>	"00001000000000110000100000000100",
		857 =>	"00000100000001000000010000000100",
		858 =>	"00000100000001000000010000000100",
		859 =>	"00000011000010110000100000001011",
		860 =>	"00001000000000110000001100000100",
		861 =>	"00000100000010110000101100001011",
		862 =>	"00001011000010110000101100000100",
		863 =>	"00000011000010110000100000001011",
		864 =>	"00001000000000110000101100000011",
		865 =>	"00000011000001000000010000001011",
		866 =>	"00000100000001000000010000000100",
		867 =>	"00000100000000110000100000001011",
		868 =>	"00001000000000110000101100001011",
		869 =>	"00001011000000110000010000000011",
		870 =>	"00000011000001000000100000001011",
		871 =>	"00000100000000110000100000001011",
		872 =>	"00001000000000110000101100001011",
		873 =>	"00001011000010110000001100000100",
		874 =>	"00000100000001000000100000001011",
		875 =>	"00000100000000110000100000001011",
		876 =>	"00001000000000110000101100001011",
		877 =>	"00001011000010110000101100000011",
		878 =>	"00000011000001000000101100001011",
		879 =>	"00000100000000110000100000001011",
		880 =>	"00001000000000110000101100001011",
		881 =>	"00001011000010110000101100001011",
		882 =>	"00001011000001000000010000000100",
		883 =>	"00000100000000110000100000001011",
		884 =>	"00001000000000110000101100001011",
		885 =>	"00001011000010110000101100001011",
		886 =>	"00001011000000110000001100000011",
		887 =>	"00000011000010110000100000001011",
		888 =>	"00000100000010000000100000001000",
		889 =>	"00001000000010000000100000001000",
		890 =>	"00001000000010000000100000001000",
		891 =>	"00001000000010000000010000001011",
		892 =>	"00000011000010110000101100001011",
		893 =>	"00001011000010110000101100001011",
		894 =>	"00001011000010110000101100001011",
		895 =>	"00001011000010110000101100000011",
		896 =>	"00000011000000110000001100000011", -- IMG_16x16_BONUS_TIME
		897 =>	"00000011000000110000001100000011",
		898 =>	"00000011000000110000001100000011",
		899 =>	"00000011000000110000001100000011",
		900 =>	"00000011000000110000100000001000",
		901 =>	"00001000000010000000100000001000",
		902 =>	"00001000000010000000100000001000",
		903 =>	"00001000000010000000100000000100",
		904 =>	"00001011000010000000001100000011",
		905 =>	"00000011000000110000001100000011",
		906 =>	"00000011000000110000001100000011",
		907 =>	"00000011000000110000001100001000",
		908 =>	"00001011000010000000001100001011",
		909 =>	"00001011000010110000101100001000",
		910 =>	"00000100000010000000010000000011",
		911 =>	"00001011000010110000101100001000",
		912 =>	"00001011000010000000001100001011",
		913 =>	"00001011000010110000101100000100",
		914 =>	"00000011000000110000001100001000",
		915 =>	"00000100000000110000101100001000",
		916 =>	"00001011000010000000001100001011",
		917 =>	"00001011000010110000010000000100",
		918 =>	"00000100000001000000001100000011",
		919 =>	"00000011000000110000101100001000",
		920 =>	"00001011000010000000001100001011",
		921 =>	"00001011000001000000100000001000",
		922 =>	"00001000000010000000010000000011",
		923 =>	"00001011000010110000101100001000",
		924 =>	"00001011000010000000001100001011",
		925 =>	"00000100000010000000100000001011",
		926 =>	"00001000000010000000100000000100",
		927 =>	"00000011000010110000101100001000",
		928 =>	"00001011000010000000001100001011",
		929 =>	"00000100000010000000100000001011",
		930 =>	"00001000000010000000100000000100",
		931 =>	"00000011000010110000101100001000",
		932 =>	"00001011000010000000001100001011",
		933 =>	"00000100000010000000100000001000",
		934 =>	"00001011000010000000100000000100",
		935 =>	"00000011000010110000101100001000",
		936 =>	"00001011000010000000001100001011",
		937 =>	"00000011000001000000100000001000",
		938 =>	"00001000000010000000010000000011",
		939 =>	"00001011000010110000101100001000",
		940 =>	"00001011000010000000001100001011",
		941 =>	"00001011000000110000010000000100",
		942 =>	"00000100000001000000001100001011",
		943 =>	"00001011000010110000101100001000",
		944 =>	"00001011000010000000001100001011",
		945 =>	"00001011000010110000001100000011",
		946 =>	"00000011000000110000101100001011",
		947 =>	"00001011000010110000101100001000",
		948 =>	"00001011000010000000001100001011",
		949 =>	"00001011000010110000101100001011",
		950 =>	"00001011000010110000101100001011",
		951 =>	"00001011000010110000101100001000",
		952 =>	"00001011000001000000100000001000",
		953 =>	"00001000000010000000100000001000",
		954 =>	"00001000000010000000100000001000",
		955 =>	"00001000000010000000100000000100",
		956 =>	"00000011000000110000101100001011",
		957 =>	"00001011000010110000101100001011",
		958 =>	"00001011000010110000101100001011",
		959 =>	"00001011000010110000101100001011",
		960 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK1
		961 =>	"00000011000000110000001100000011",
		962 =>	"00000011000000110000001100000011",
		963 =>	"00000011000000110000001100000011",
		964 =>	"00000011000000110000001100000011",
		965 =>	"00000011000000110000001100001000",
		966 =>	"00000011000000110000001100000011",
		967 =>	"00000011000000110000001100000011",
		968 =>	"00000011000000110000001100000011",
		969 =>	"00000011000000110000001100001000",
		970 =>	"00000011000000110000001100000011",
		971 =>	"00000011000000110000001100000011",
		972 =>	"00000011000000110000001100000011",
		973 =>	"00000011000000110000001100001000",
		974 =>	"00000011000000110000001100000011",
		975 =>	"00000011000000110000001100000011",
		976 =>	"00000011000010000000010000000100",
		977 =>	"00000011000000110000010000001000",
		978 =>	"00001011000000110000001100001000",
		979 =>	"00000100000001000000001100000011",
		980 =>	"00000011000010110000101100000100",
		981 =>	"00000011000010000000010000001000",
		982 =>	"00001011000010110000001100000100",
		983 =>	"00001011000010110000001100000011",
		984 =>	"00000011000010000000010000000100",
		985 =>	"00001000000010000000010000001000",
		986 =>	"00001011000010110000101100000100",
		987 =>	"00000100000001000000001100000011",
		988 =>	"00000011000010110000101100000100",
		989 =>	"00001000000010000000010000000100",
		990 =>	"00000100000010110000101100000100",
		991 =>	"00001011000010110000001100000011",
		992 =>	"00000011000010000000010000000100",
		993 =>	"00001000000001000000010000001011",
		994 =>	"00000100000001000000101100000100",
		995 =>	"00000100000001000000001100000011",
		996 =>	"00000011000010110000101100000100",
		997 =>	"00001000000001000000101100001011",
		998 =>	"00001000000001000000101100000100",
		999 =>	"00001011000010110000001100000011",
		1000 =>	"00000011000010000000010000000100",
		1001 =>	"00001000000001000000101100001000",
		1002 =>	"00001000000001000000101100000100",
		1003 =>	"00000100000001000000001100000011",
		1004 =>	"00000011000010110000101100000100",
		1005 =>	"00001000000001000000010000000100",
		1006 =>	"00000100000001000000101100000100",
		1007 =>	"00001011000010110000001100000011",
		1008 =>	"00000011000010000000010000000100",
		1009 =>	"00001000000010000000010000000100",
		1010 =>	"00000100000010110000101100000100",
		1011 =>	"00000100000001000000001100000011",
		1012 =>	"00000011000010110000101100000100",
		1013 =>	"00000011000010000000010000000100",
		1014 =>	"00001011000010110000001100000100",
		1015 =>	"00001011000010110000001100000011",
		1016 =>	"00000011000010000000010000000100",
		1017 =>	"00000011000000110000101100001011",
		1018 =>	"00001011000000110000001100000100",
		1019 =>	"00000100000001000000001100000011",
		1020 =>	"00000011000000110000001100000011",
		1021 =>	"00000011000000110000001100000100",
		1022 =>	"00000011000000110000001100000011",
		1023 =>	"00000011000000110000001100000011",
		1024 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK2
		1025 =>	"00000011000000110000001100000011",
		1026 =>	"00000011000000110000001100000011",
		1027 =>	"00000011000000110000001100000011",
		1028 =>	"00000011000000110000001100000011",
		1029 =>	"00000011000000110000001100001000",
		1030 =>	"00000011000000110000001100000011",
		1031 =>	"00000011000000110000001100000011",
		1032 =>	"00000011000000110000001100000011",
		1033 =>	"00000011000000110000001100001000",
		1034 =>	"00000011000000110000001100000011",
		1035 =>	"00000011000000110000001100000011",
		1036 =>	"00000011000001000000101100000011",
		1037 =>	"00001000000010000000101100001000",
		1038 =>	"00001011000001000000010000000011",
		1039 =>	"00000100000010110000001100000011",
		1040 =>	"00000011000010110000101100001000",
		1041 =>	"00001000000010000000101100001000",
		1042 =>	"00001011000001000000010000000100",
		1043 =>	"00001011000010110000001100000011",
		1044 =>	"00000011000010110000101100000100",
		1045 =>	"00001000000010000000101100001000",
		1046 =>	"00001011000010110000101100000100",
		1047 =>	"00001011000010110000001100000011",
		1048 =>	"00000011000000110000001100000100",
		1049 =>	"00000100000010000000010000001000",
		1050 =>	"00000100000010110000101100000100",
		1051 =>	"00000011000000110000001100000011",
		1052 =>	"00000011000000110000001100000100",
		1053 =>	"00001000000001000000010000000100",
		1054 =>	"00000100000001000000101100000100",
		1055 =>	"00000011000000110000001100000011",
		1056 =>	"00000011000001000000101100000100",
		1057 =>	"00001000000001000000010000001011",
		1058 =>	"00000100000001000000101100000100",
		1059 =>	"00000100000010110000001100000011",
		1060 =>	"00000011000010110000101100000100",
		1061 =>	"00001000000001000000101100001011",
		1062 =>	"00001000000001000000101100000100",
		1063 =>	"00001011000010110000001100000011",
		1064 =>	"00000011000010110000101100000100",
		1065 =>	"00001000000001000000101100001000",
		1066 =>	"00001000000001000000101100000100",
		1067 =>	"00001011000010110000001100000011",
		1068 =>	"00000011000000110000001100000100",
		1069 =>	"00001000000001000000010000000100",
		1070 =>	"00000100000001000000101100000100",
		1071 =>	"00000011000000110000001100000011",
		1072 =>	"00000011000000110000001100000100",
		1073 =>	"00001000000010000000010000000100",
		1074 =>	"00000100000010000000101100000100",
		1075 =>	"00000011000000110000001100000011",
		1076 =>	"00000011000001000000101100000100",
		1077 =>	"00000100000001000000100000001000",
		1078 =>	"00001000000010110000101100000100",
		1079 =>	"00000100000010110000001100000011",
		1080 =>	"00000011000010110000101100000100",
		1081 =>	"00001011000010110000101100001011",
		1082 =>	"00001011000010110000101100000100",
		1083 =>	"00001011000010110000001100000011",
		1084 =>	"00000011000010110000101100000011",
		1085 =>	"00001011000010110000101100001000",
		1086 =>	"00001011000010110000101100000011",
		1087 =>	"00001011000010110000001100000011",
		1088 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK3
		1089 =>	"00000011000000110000001100000011",
		1090 =>	"00000011000000110000001100000011",
		1091 =>	"00000011000000110000001100000011",
		1092 =>	"00000011000000110000001100000011",
		1093 =>	"00000011000000110000100000001000",
		1094 =>	"00000100000000110000001100000011",
		1095 =>	"00000011000000110000001100000011",
		1096 =>	"00000011000000110000001100000011",
		1097 =>	"00000011000000110000001100001000",
		1098 =>	"00000011000000110000001100000011",
		1099 =>	"00000011000000110000001100000011",
		1100 =>	"00000011000000110000001100000011",
		1101 =>	"00000011000000110000001100001000",
		1102 =>	"00000011000000110000001100000011",
		1103 =>	"00000011000000110000001100000011",
		1104 =>	"00000011000010000000010000000100",
		1105 =>	"00000011000000110000010000001000",
		1106 =>	"00001011000000110000001100001000",
		1107 =>	"00000100000001000000001100000011",
		1108 =>	"00000011000010110000101100000100",
		1109 =>	"00000011000010000000010000001000",
		1110 =>	"00001011000010110000001100000100",
		1111 =>	"00001011000010110000001100000011",
		1112 =>	"00000011000010000000010000000100",
		1113 =>	"00001000000010000000010000001000",
		1114 =>	"00001011000010110000101100000100",
		1115 =>	"00000100000001000000001100000011",
		1116 =>	"00000011000010110000101100000100",
		1117 =>	"00001000000010000000010000000100",
		1118 =>	"00000100000010110000101100000100",
		1119 =>	"00001011000010110000001100000011",
		1120 =>	"00000011000010000000010000000100",
		1121 =>	"00001000000001000000010000001011",
		1122 =>	"00000100000001000000101100000100",
		1123 =>	"00000100000001000000001100000011",
		1124 =>	"00000011000010110000101100000100",
		1125 =>	"00001000000001000000101100001011",
		1126 =>	"00001000000001000000101100000100",
		1127 =>	"00001011000010110000001100000011",
		1128 =>	"00000011000010000000010000000100",
		1129 =>	"00001000000001000000101100001000",
		1130 =>	"00001000000001000000101100000100",
		1131 =>	"00000100000001000000001100000011",
		1132 =>	"00000011000010110000101100000100",
		1133 =>	"00001000000001000000010000000100",
		1134 =>	"00000100000001000000101100000100",
		1135 =>	"00001011000010110000001100000011",
		1136 =>	"00000011000010000000010000000100",
		1137 =>	"00001000000010000000010000000100",
		1138 =>	"00000100000010110000101100000100",
		1139 =>	"00000100000001000000001100000011",
		1140 =>	"00000011000010110000101100000100",
		1141 =>	"00000011000010000000100000000100",
		1142 =>	"00001011000010110000001100000100",
		1143 =>	"00001011000010110000001100000011",
		1144 =>	"00000011000010000000010000000100",
		1145 =>	"00000011000010000000100000001011",
		1146 =>	"00001011000010110000001100000100",
		1147 =>	"00000100000001000000001100000011",
		1148 =>	"00000011000010110000101100000100",
		1149 =>	"00000011000000110000010000001000",
		1150 =>	"00001011000000110000001100000100",
		1151 =>	"00001011000010110000001100000011",
		1152 =>	"00000011000000110000001100000011", -- IMG_16x16_ENEMY_TANK4
		1153 =>	"00000011000000110000001100000011",
		1154 =>	"00000011000000110000001100000011",
		1155 =>	"00000011000000110000001100000011",
		1156 =>	"00000011000010000000010000000100",
		1157 =>	"00000011000000110000100000001000",
		1158 =>	"00000100000000110000001100001000",
		1159 =>	"00000100000001000000001100000011",
		1160 =>	"00000011000010110000101100000100",
		1161 =>	"00000100000010110000100000001000",
		1162 =>	"00000100000010110000010000000100",
		1163 =>	"00001011000010110000001100000011",
		1164 =>	"00000011000010000000010000000100",
		1165 =>	"00000100000001000000010000001000",
		1166 =>	"00001011000001000000010000000100",
		1167 =>	"00000100000001000000001100000011",
		1168 =>	"00000011000010110000101100000100",
		1169 =>	"00001000000001000000010000001000",
		1170 =>	"00001011000001000000010000001011",
		1171 =>	"00001011000010110000001100000011",
		1172 =>	"00000011000010000000010000000100",
		1173 =>	"00001000000001000000010000001000",
		1174 =>	"00001011000010000000010000001011",
		1175 =>	"00000100000001000000001100000011",
		1176 =>	"00000011000010110000101100000100",
		1177 =>	"00001000000010000000010000001000",
		1178 =>	"00001011000010000000101100001011",
		1179 =>	"00001011000010110000001100000011",
		1180 =>	"00000011000010000000010000000100",
		1181 =>	"00001000000010000000100000001000",
		1182 =>	"00001000000010000000101100001011",
		1183 =>	"00000100000001000000001100000011",
		1184 =>	"00000011000010110000101100000100",
		1185 =>	"00001000000001000000010000001011",
		1186 =>	"00000100000001000000101100001011",
		1187 =>	"00001011000010110000001100000011",
		1188 =>	"00000011000010000000010000000100",
		1189 =>	"00001000000001000000101100001011",
		1190 =>	"00001000000001000000101100001011",
		1191 =>	"00000100000001000000001100000011",
		1192 =>	"00000011000010110000101100000100",
		1193 =>	"00001000000001000000101100001000",
		1194 =>	"00001000000001000000101100001011",
		1195 =>	"00001011000010110000001100000011",
		1196 =>	"00000011000010000000010000000100",
		1197 =>	"00001000000001000000010000000100",
		1198 =>	"00000100000001000000101100001011",
		1199 =>	"00000100000001000000001100000011",
		1200 =>	"00000011000010110000101100000100",
		1201 =>	"00001000000001000000010000000100",
		1202 =>	"00000100000001000000101100001011",
		1203 =>	"00001011000010110000001100000011",
		1204 =>	"00000011000010000000010000000100",
		1205 =>	"00000100000010110000101100001011",
		1206 =>	"00001011000010110000010000001011",
		1207 =>	"00000100000001000000001100000011",
		1208 =>	"00000011000010110000101100000100",
		1209 =>	"00001011000010110000101100001011",
		1210 =>	"00001011000010110000101100000100",
		1211 =>	"00001011000010110000001100000011",
		1212 =>	"00000011000010000000010000000100",
		1213 =>	"00000011000000110000001100000100",
		1214 =>	"00000011000000110000001100001011",
		1215 =>	"00000100000001000000001100000011",
		1216 =>	"00000011000000110000001100000011", -- IMG_16x16_EXPLOSION
		1217 =>	"00001100000000110000110000000011",
		1218 =>	"00000011000000110000001100001100",
		1219 =>	"00000011000000110000110000000011",
		1220 =>	"00000011000010000000001100000011",
		1221 =>	"00000011000010000000001100000011",
		1222 =>	"00001000000000110000110000000011",
		1223 =>	"00000011000010000000110000000011",
		1224 =>	"00000011000011000000110000001000",
		1225 =>	"00001000000000110000001100001000",
		1226 =>	"00001000000000110000001100000011",
		1227 =>	"00001000000011000000001100000011",
		1228 =>	"00000011000000110000110000001100",
		1229 =>	"00001000000011000000110000001000",
		1230 =>	"00001100000011000000001100001000",
		1231 =>	"00001000000011000000001100000011",
		1232 =>	"00000011000000110000001100001100",
		1233 =>	"00001101000010000000100000001000",
		1234 =>	"00001000000011000000100000001000",
		1235 =>	"00001100000011000000001100001100",
		1236 =>	"00000011000010000000001100001100",
		1237 =>	"00001000000010000000110100001000",
		1238 =>	"00000011000010000000100000001101",
		1239 =>	"00001100000000110000001100000011",
		1240 =>	"00000011000000110000110000001000",
		1241 =>	"00001000000011010000110000001101",
		1242 =>	"00001101000000110000110100001100",
		1243 =>	"00001000000011000000001100000011",
		1244 =>	"00001000000010000000100000001000",
		1245 =>	"00000011000010000000110100000011",
		1246 =>	"00000011000011010000100000001000",
		1247 =>	"00001000000010000000100000001000",
		1248 =>	"00000011000011000000110000001100",
		1249 =>	"00001000000010000000110000001101",
		1250 =>	"00000011000011010000100000001100",
		1251 =>	"00001100000011000000001100000011",
		1252 =>	"00000011000000110000001100001100",
		1253 =>	"00001100000011000000001100001000",
		1254 =>	"00001101000000110000110000001100",
		1255 =>	"00001000000010000000001100000011",
		1256 =>	"00000011000010000000110000001100",
		1257 =>	"00001000000010000000110000001000",
		1258 =>	"00000011000010000000110100001000",
		1259 =>	"00001100000011000000100000000011",
		1260 =>	"00000011000000110000100000001000",
		1261 =>	"00001000000011010000100000001100",
		1262 =>	"00001000000011000000100000001000",
		1263 =>	"00000011000000110000001100000011",
		1264 =>	"00000011000011000000100000001100",
		1265 =>	"00001100000010000000110000001000",
		1266 =>	"00001000000011000000110000001000",
		1267 =>	"00001000000000110000110000000011",
		1268 =>	"00000011000010000000110000000011",
		1269 =>	"00000011000011000000001100001100",
		1270 =>	"00001000000011000000001100001100",
		1271 =>	"00001100000010000000001100000011",
		1272 =>	"00001000000011000000001100000011",
		1273 =>	"00001100000000110000001100000011",
		1274 =>	"00001000000000110000001100000011",
		1275 =>	"00000011000011000000100000000011",
		1276 =>	"00000011000000110000001100000011",
		1277 =>	"00000011000000110000001100000011",
		1278 =>	"00001000000000110000110000000011",
		1279 =>	"00000011000000110000110000000011",
		1280 =>	"00000011000000110000000100000001", -- IMG_16x16_FLAG
		1281 =>	"00000001000000010000000100000001",
		1282 =>	"00000001000000010000000100000001",
		1283 =>	"00000001000000010000000100000001",
		1284 =>	"00000011000000110000001000000010",
		1285 =>	"00000001000000010000000100000001",
		1286 =>	"00000001000000010000000100000001",
		1287 =>	"00000001000000010000000100000001",
		1288 =>	"00000011000000110000001000000010",
		1289 =>	"00000010000000100000000100000001",
		1290 =>	"00000001000000010000000100000001",
		1291 =>	"00000001000000010000000100000001",
		1292 =>	"00000011000000110000001000000010",
		1293 =>	"00000010000000100000001000000010",
		1294 =>	"00000001000000010000000100000001",
		1295 =>	"00000001000000010000000100000001",
		1296 =>	"00000011000000110000001000000010",
		1297 =>	"00000010000000100000001000000010",
		1298 =>	"00000010000000100000000100000001",
		1299 =>	"00000001000000010000000100000001",
		1300 =>	"00000011000000110000001000000010",
		1301 =>	"00000010000000100000001000000010",
		1302 =>	"00000010000000100000001000000010",
		1303 =>	"00000001000000010000000100000001",
		1304 =>	"00000011000000110000001000000010",
		1305 =>	"00000010000000100000001000000010",
		1306 =>	"00000010000000100000001000000010",
		1307 =>	"00000010000000100000000100000001",
		1308 =>	"00000011000000110000001000000010",
		1309 =>	"00000010000000100000001000000010",
		1310 =>	"00000010000000100000001000000010",
		1311 =>	"00000010000000100000001000000010",
		1312 =>	"00000011000000110000001000000010",
		1313 =>	"00000010000000100000001000000010",
		1314 =>	"00000010000000100000001000000010",
		1315 =>	"00000010000000100000001000000010",
		1316 =>	"00000011000000110000000100000001",
		1317 =>	"00000001000000010000000100000001",
		1318 =>	"00000001000000010000000100000001",
		1319 =>	"00000001000000010000000100000001",
		1320 =>	"00000011000000110000000100000001",
		1321 =>	"00000001000000010000000100000001",
		1322 =>	"00000001000000010000000100000001",
		1323 =>	"00000001000000010000000100000001",
		1324 =>	"00000011000000110000000100000001",
		1325 =>	"00000001000000010000000100000001",
		1326 =>	"00000001000000010000000100000001",
		1327 =>	"00000001000000010000000100000001",
		1328 =>	"00000011000000110000000100000001",
		1329 =>	"00000001000000010000000100000001",
		1330 =>	"00000001000000010000000100000001",
		1331 =>	"00000001000000010000000100000001",
		1332 =>	"00000011000000110000000100000001",
		1333 =>	"00000001000000010000000100000001",
		1334 =>	"00000001000000010000000100000001",
		1335 =>	"00000001000000010000000100000001",
		1336 =>	"00000011000000110000000100000001",
		1337 =>	"00000001000000010000000100000001",
		1338 =>	"00000001000000010000000100000001",
		1339 =>	"00000001000000010000000100000001",
		1340 =>	"00000001000000010000000100000001",
		1341 =>	"00000001000000010000000100000001",
		1342 =>	"00000001000000010000000100000001",
		1343 =>	"00000001000000010000000100000001",
		1344 =>	"00000011000000110000001100000011", -- IMG_16x16_MAIN_TANK
		1345 =>	"00000011000000110000001100000011",
		1346 =>	"00000011000000110000001100000011",
		1347 =>	"00000011000000110000001100000011",
		1348 =>	"00000011000000110000001100000011",
		1349 =>	"00000011000000110000001100000011",
		1350 =>	"00000011000000110000001100000011",
		1351 =>	"00000011000000110000001100000011",
		1352 =>	"00000011000000110000001100000011",
		1353 =>	"00000011000000110000001100001110",
		1354 =>	"00000011000000110000001100000011",
		1355 =>	"00000011000000110000001100000011",
		1356 =>	"00000011000000110000001100000011",
		1357 =>	"00000011000000110000001100001110",
		1358 =>	"00000011000000110000001100000011",
		1359 =>	"00000011000000110000001100000011",
		1360 =>	"00000011000011100000111100001111",
		1361 =>	"00000011000000110000001100001110",
		1362 =>	"00000011000000110000001100001110",
		1363 =>	"00001111000011110000001100000011",
		1364 =>	"00000011000100000001000000001110",
		1365 =>	"00000011000000110000001100001110",
		1366 =>	"00000011000000110000001100010000",
		1367 =>	"00010000000100000000001100000011",
		1368 =>	"00000011000011100000111100001110",
		1369 =>	"00000011000011100000111100001110",
		1370 =>	"00010000000100000000001100010000",
		1371 =>	"00001111000011110000001100000011",
		1372 =>	"00000011000100000001000000001110",
		1373 =>	"00001110000011100000111100001111",
		1374 =>	"00001111000011110001000000010000",
		1375 =>	"00010000000100000000001100000011",
		1376 =>	"00000011000011100000111100001110",
		1377 =>	"00001110000011110000111000001110",
		1378 =>	"00001111000011110000111100010000",
		1379 =>	"00001111000011110000001100000011",
		1380 =>	"00000011000100000001000000001110",
		1381 =>	"00001110000011110000111000001111",
		1382 =>	"00010000000011110000111100010000",
		1383 =>	"00010000000100000000001100000011",
		1384 =>	"00000011000011100000111100001110",
		1385 =>	"00001110000011110000111000001111",
		1386 =>	"00010000000011110000111100010000",
		1387 =>	"00001111000011110000001100000011",
		1388 =>	"00000011000100000001000000001110",
		1389 =>	"00001110000011100000111100010000",
		1390 =>	"00010000000011110000111100010000",
		1391 =>	"00010000000100000000001100000011",
		1392 =>	"00000011000011100000111100001110",
		1393 =>	"00010000000011100000111000001111",
		1394 =>	"00001111000011110001000000010000",
		1395 =>	"00001111000011110000001100000011",
		1396 =>	"00000011000100000001000000001110",
		1397 =>	"00000011000100000001000000010000",
		1398 =>	"00010000000100000000001100010000",
		1399 =>	"00010000000100000000001100000011",
		1400 =>	"00000011000011100000111100001111",
		1401 =>	"00000011000000110000001100000011",
		1402 =>	"00000011000000110000001100010000",
		1403 =>	"00001111000011110000001100000011",
		1404 =>	"00000011000000110000001100000011",
		1405 =>	"00000011000000110000001100000011",
		1406 =>	"00000011000000110000001100000011",
		1407 =>	"00000011000000110000001100000011",


--			***** MAP *****


		1408 =>	"00000010000000000000000100000000", -- z: 2 rot: 0 ptr: 256
		1409 =>	"00000010000000000000000100010000", -- z: 2 rot: 0 ptr: 272
		1410 =>	"00000011000000000000000100100000", -- z: 3 rot: 0 ptr: 288
		1411 =>	"00000001000000000000000100110000", -- z: 1 rot: 0 ptr: 304
		1412 =>	"00000010000000000000000101000000", -- z: 2 rot: 0 ptr: 320
		1413 =>	"00000010000000000000000101010000", -- z: 2 rot: 0 ptr: 336
		1414 =>	"00000010000000000000000101100000", -- z: 2 rot: 0 ptr: 352
		1415 =>	"00000001000000000000000101110000", -- z: 1 rot: 0 ptr: 368
		1416 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1417 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1418 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1419 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1420 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1421 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1422 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1423 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1424 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1425 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1426 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1427 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1428 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1429 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1430 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1431 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1432 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1433 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1434 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1435 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1436 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1437 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1438 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1439 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1440 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1441 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1442 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1443 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1444 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1445 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1446 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1447 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1448 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1449 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1450 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1451 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1452 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1453 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1454 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1455 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1456 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1457 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1458 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1459 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1460 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1461 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1462 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1463 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1464 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1465 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1466 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1467 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1468 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1469 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1470 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1471 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1472 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1473 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1474 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1475 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1476 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1477 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1478 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1479 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1480 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1481 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1482 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1483 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1484 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1485 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1486 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1487 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1488 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1489 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1490 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1491 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1492 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1493 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1494 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1495 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1496 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1497 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1498 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1499 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1500 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1501 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1502 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1503 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1504 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1505 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1506 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1507 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1508 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1509 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1510 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1511 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1512 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1513 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1514 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1515 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1516 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1517 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1518 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1519 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1520 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1521 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1522 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1523 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1524 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1525 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1526 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1527 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1528 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1529 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1530 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1531 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1532 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1533 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1534 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1535 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1536 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1537 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1538 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1539 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1540 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1541 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1542 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1543 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1544 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1545 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1546 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1547 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1548 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1549 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1550 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1551 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1552 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1553 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1554 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1555 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1556 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1557 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1558 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1559 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1560 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1561 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1562 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1563 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1564 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1565 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1566 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1567 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1568 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1569 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1570 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1571 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1572 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1573 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1574 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1575 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1576 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1577 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1578 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1579 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1580 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1581 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1582 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1583 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1584 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1585 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1586 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1587 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1588 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1589 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1590 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1591 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1592 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1593 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1594 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1595 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1596 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1597 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1598 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1599 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1600 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1601 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1602 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1603 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1604 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1605 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1606 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1607 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1608 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1609 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1610 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1611 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1612 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1613 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1614 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1615 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1616 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1617 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1618 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1619 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1620 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1621 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1622 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1623 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1624 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1625 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1626 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1627 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1628 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1629 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1630 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1631 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1632 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1633 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1634 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1635 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1636 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1637 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1638 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1639 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1640 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1641 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1642 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1643 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1644 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1645 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1646 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1647 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1648 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1649 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1650 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1651 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1652 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1653 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1654 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1655 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1656 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1657 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1658 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1659 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1660 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1661 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1662 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1663 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1664 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1665 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1666 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1667 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1668 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1669 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1670 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1671 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1672 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1673 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1674 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1675 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1676 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1677 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1678 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1679 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1680 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1681 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1682 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1683 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1684 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1685 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1686 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1687 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1688 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1689 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1690 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1691 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1692 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1693 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1694 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1695 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1696 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1697 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1698 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1699 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1700 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1701 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1702 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1703 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1704 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1705 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1706 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1707 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1708 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1709 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1710 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1711 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1712 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1713 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1714 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1715 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1716 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1717 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1718 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1719 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1720 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1721 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1722 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1723 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1724 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1725 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1726 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1727 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1728 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1729 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1730 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1731 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1732 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1733 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1734 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1735 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1736 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1737 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1738 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1739 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1740 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1741 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1742 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1743 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1744 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1745 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1746 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1747 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1748 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1749 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1750 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1751 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1752 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1753 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1754 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1755 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1756 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1757 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1758 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1759 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1760 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1761 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1762 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1763 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1764 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1765 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1766 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1767 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1768 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1769 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1770 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1771 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1772 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1773 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1774 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1775 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1776 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1777 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1778 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1779 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1780 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1781 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1782 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1783 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1784 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1785 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1786 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1787 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1788 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1789 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1790 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1791 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1792 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1793 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1794 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1795 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1796 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1797 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1798 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1799 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1800 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1801 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1802 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1803 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1804 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1805 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1806 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1807 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1808 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1809 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1810 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1811 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1812 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1813 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1814 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1815 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1816 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1817 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1818 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1819 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1820 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1821 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1822 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1823 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1824 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1825 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1826 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1827 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1828 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1829 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1830 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1831 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1832 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1833 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1834 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1835 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1836 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1837 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1838 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1839 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1840 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1841 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1842 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1843 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1844 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1845 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1846 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1847 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1848 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1849 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1850 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1851 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1852 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1853 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1854 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1855 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1856 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1857 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1858 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1859 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1860 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1861 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1862 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1863 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1864 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1865 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1866 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1867 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1868 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1869 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1870 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1871 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1872 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1873 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1874 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1875 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1876 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1877 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1878 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1879 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1880 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1881 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1882 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1883 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1884 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1885 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1886 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1887 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1888 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1889 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1890 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1891 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1892 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1893 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1894 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1895 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1896 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1897 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1898 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1899 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1900 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1901 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1902 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1903 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1904 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1905 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1906 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1907 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1908 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1909 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1910 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1911 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1912 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1913 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1914 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1915 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1916 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1917 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1918 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1919 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1920 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1921 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1922 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1923 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1924 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1925 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1926 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1927 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1928 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1929 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1930 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1931 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1932 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1933 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1934 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1935 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1936 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1937 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1938 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1939 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1940 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1941 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1942 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1943 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1944 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1945 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1946 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1947 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1948 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1949 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1950 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1951 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1952 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1953 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1954 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1955 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1956 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1957 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1958 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1959 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1960 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1961 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1962 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1963 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1964 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1965 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1966 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1967 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1968 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1969 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1970 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1971 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1972 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1973 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1974 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1975 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1976 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1977 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1978 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1979 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1980 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1981 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1982 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1983 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1984 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1985 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1986 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1987 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1988 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1989 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1990 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1991 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1992 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1993 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1994 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1995 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1996 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1997 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1998 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		1999 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2000 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2001 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2002 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2003 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2004 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2005 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2006 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2007 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2008 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2009 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2010 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2011 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2012 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2013 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2014 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2015 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2016 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2017 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2018 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2019 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2020 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2021 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2022 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2023 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2024 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2025 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2026 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2027 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2028 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2029 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2030 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2031 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2032 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2033 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2034 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2035 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2036 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2037 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2038 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2039 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2040 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2041 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2042 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2043 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2044 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2045 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2046 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2047 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2048 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2049 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2050 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2051 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2052 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2053 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2054 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2055 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2056 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2057 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2058 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2059 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2060 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2061 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2062 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2063 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2064 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2065 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2066 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2067 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2068 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2069 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2070 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2071 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2072 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2073 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2074 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2075 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2076 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2077 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2078 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2079 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2080 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2081 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2082 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2083 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2084 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2085 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2086 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2087 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2088 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2089 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2090 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2091 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2092 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2093 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2094 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2095 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2096 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2097 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2098 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2099 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2100 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2101 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2102 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2103 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2104 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2105 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2106 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2107 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2108 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2109 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2110 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2111 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2112 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2113 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2114 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2115 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2116 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2117 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2118 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2119 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2120 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2121 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2122 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2123 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2124 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2125 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2126 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2127 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2128 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2129 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2130 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2131 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2132 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2133 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2134 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2135 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2136 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2137 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2138 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2139 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2140 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2141 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2142 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2143 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2144 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2145 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2146 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2147 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2148 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2149 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2150 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2151 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2152 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2153 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2154 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2155 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2156 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2157 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2158 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2159 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2160 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2161 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2162 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2163 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2164 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2165 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2166 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2167 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2168 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2169 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2170 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2171 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2172 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2173 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2174 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2175 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2176 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2177 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2178 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2179 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2180 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2181 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2182 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2183 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2184 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2185 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2186 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2187 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2188 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2189 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2190 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2191 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2192 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2193 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2194 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2195 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2196 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2197 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2198 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2199 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2200 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2201 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2202 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2203 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2204 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2205 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2206 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2207 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2208 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2209 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2210 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2211 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2212 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2213 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2214 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2215 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2216 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2217 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2218 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2219 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2220 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2221 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2222 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2223 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2224 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2225 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2226 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2227 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2228 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2229 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2230 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2231 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2232 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2233 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2234 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2235 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2236 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2237 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2238 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2239 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2240 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2241 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2242 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2243 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2244 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2245 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2246 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2247 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2248 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2249 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2250 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2251 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2252 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2253 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2254 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2255 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2256 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2257 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2258 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2259 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2260 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2261 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2262 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2263 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2264 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2265 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2266 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2267 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2268 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2269 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2270 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2271 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2272 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2273 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2274 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2275 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2276 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2277 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2278 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2279 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2280 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2281 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2282 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2283 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2284 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2285 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2286 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2287 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2288 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2289 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2290 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2291 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2292 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2293 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2294 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2295 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2296 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2297 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2298 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2299 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2300 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2301 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2302 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2303 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2304 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2305 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2306 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2307 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2308 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2309 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2310 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2311 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2312 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2313 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2314 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2315 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2316 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2317 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2318 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2319 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2320 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2321 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2322 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2323 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2324 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2325 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2326 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2327 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2328 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2329 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2330 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2331 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2332 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2333 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2334 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2335 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2336 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2337 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2338 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2339 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2340 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2341 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2342 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2343 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2344 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2345 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2346 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2347 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2348 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2349 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2350 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2351 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2352 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2353 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2354 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2355 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2356 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2357 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2358 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2359 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2360 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2361 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2362 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2363 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2364 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2365 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2366 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2367 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2368 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2369 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2370 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2371 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2372 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2373 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2374 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2375 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2376 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2377 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2378 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2379 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2380 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2381 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2382 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2383 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2384 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2385 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2386 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2387 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2388 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2389 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2390 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2391 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2392 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2393 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2394 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2395 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2396 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2397 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2398 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2399 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2400 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2401 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2402 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2403 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2404 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2405 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2406 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2407 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2408 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2409 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2410 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2411 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2412 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2413 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2414 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2415 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2416 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2417 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2418 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2419 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2420 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2421 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2422 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2423 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2424 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2425 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2426 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2427 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2428 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2429 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2430 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2431 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2432 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2433 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2434 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2435 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2436 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2437 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2438 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2439 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2440 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2441 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2442 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2443 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2444 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2445 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2446 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2447 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2448 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2449 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2450 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2451 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2452 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2453 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2454 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2455 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2456 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2457 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2458 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2459 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2460 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2461 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2462 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2463 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2464 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2465 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2466 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2467 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2468 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2469 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2470 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2471 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2472 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2473 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2474 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2475 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2476 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2477 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2478 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2479 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2480 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2481 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2482 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2483 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2484 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2485 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2486 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2487 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2488 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2489 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2490 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2491 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2492 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2493 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2494 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2495 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2496 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2497 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2498 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2499 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2500 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2501 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2502 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2503 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2504 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2505 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2506 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2507 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2508 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2509 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2510 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2511 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2512 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2513 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2514 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2515 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2516 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2517 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2518 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2519 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2520 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2521 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2522 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2523 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2524 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2525 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2526 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2527 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2528 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2529 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2530 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2531 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2532 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2533 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2534 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2535 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2536 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2537 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2538 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2539 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2540 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2541 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2542 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2543 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2544 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2545 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2546 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2547 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2548 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2549 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2550 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2551 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2552 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2553 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2554 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2555 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2556 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2557 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2558 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2559 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2560 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2561 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2562 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2563 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2564 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2565 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2566 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2567 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2568 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2569 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2570 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2571 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2572 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2573 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2574 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2575 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2576 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2577 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2578 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2579 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2580 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2581 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2582 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2583 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2584 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2585 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2586 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2587 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2588 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2589 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2590 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2591 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2592 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2593 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2594 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2595 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2596 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2597 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2598 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2599 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2600 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2601 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2602 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2603 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2604 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2605 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2606 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2607 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2608 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2609 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2610 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2611 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2612 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2613 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2614 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2615 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2616 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2617 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2618 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2619 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2620 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2621 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2622 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2623 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2624 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2625 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2626 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2627 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2628 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2629 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2630 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2631 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2632 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2633 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2634 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2635 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2636 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2637 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2638 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2639 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2640 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2641 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2642 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2643 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2644 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2645 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2646 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2647 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2648 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2649 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2650 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2651 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2652 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2653 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2654 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2655 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2656 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2657 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2658 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2659 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2660 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2661 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2662 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2663 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2664 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2665 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2666 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2667 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2668 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2669 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2670 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2671 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2672 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2673 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2674 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2675 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2676 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2677 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2678 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2679 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2680 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2681 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2682 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2683 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2684 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2685 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2686 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2687 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2688 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2689 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2690 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2691 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2692 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2693 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2694 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2695 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2696 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2697 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2698 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2699 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2700 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2701 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2702 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2703 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2704 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2705 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2706 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2707 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2708 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2709 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2710 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2711 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2712 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2713 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2714 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2715 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2716 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2717 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2718 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2719 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2720 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2721 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2722 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2723 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2724 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2725 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2726 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2727 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2728 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2729 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2730 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2731 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2732 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2733 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2734 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2735 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2736 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2737 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2738 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2739 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2740 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2741 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2742 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2743 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2744 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2745 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2746 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2747 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2748 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2749 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2750 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2751 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2752 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2753 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2754 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2755 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2756 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2757 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2758 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2759 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2760 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2761 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2762 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2763 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2764 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2765 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2766 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2767 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2768 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2769 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2770 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2771 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2772 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2773 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2774 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2775 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2776 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2777 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2778 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2779 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2780 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2781 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2782 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2783 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2784 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2785 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2786 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2787 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2788 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2789 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2790 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2791 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2792 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2793 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2794 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2795 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2796 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2797 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2798 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2799 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2800 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2801 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2802 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2803 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2804 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2805 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2806 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2807 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2808 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2809 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2810 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2811 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2812 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2813 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2814 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2815 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2816 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2817 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2818 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2819 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2820 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2821 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2822 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2823 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2824 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2825 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2826 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2827 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2828 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2829 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2830 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2831 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2832 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2833 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2834 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2835 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2836 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2837 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2838 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2839 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2840 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2841 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2842 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2843 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2844 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2845 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2846 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2847 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2848 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2849 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2850 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2851 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2852 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2853 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2854 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2855 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2856 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2857 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2858 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2859 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2860 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2861 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2862 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2863 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2864 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2865 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2866 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2867 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2868 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2869 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2870 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2871 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2872 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2873 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2874 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2875 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2876 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2877 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2878 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2879 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2880 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2881 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2882 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2883 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2884 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2885 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2886 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2887 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2888 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2889 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2890 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2891 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2892 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2893 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2894 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2895 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2896 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2897 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2898 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2899 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2900 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2901 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2902 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2903 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2904 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2905 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2906 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2907 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2908 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2909 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2910 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2911 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2912 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2913 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2914 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2915 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2916 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2917 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2918 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2919 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2920 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2921 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2922 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2923 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2924 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2925 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2926 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2927 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2928 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2929 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2930 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2931 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2932 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2933 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2934 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2935 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2936 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2937 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2938 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2939 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2940 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2941 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2942 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2943 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2944 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2945 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2946 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2947 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2948 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2949 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2950 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2951 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2952 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2953 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2954 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2955 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2956 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2957 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2958 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2959 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2960 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2961 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2962 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2963 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2964 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2965 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2966 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2967 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2968 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2969 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2970 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2971 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2972 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2973 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2974 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2975 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2976 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2977 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2978 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2979 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2980 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2981 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2982 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2983 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2984 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2985 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2986 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2987 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2988 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2989 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2990 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2991 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2992 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2993 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2994 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2995 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2996 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2997 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2998 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		2999 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3000 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3001 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3002 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3003 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3004 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3005 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3006 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3007 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3008 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3009 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3010 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3011 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3012 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3013 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3014 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3015 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3016 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3017 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3018 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3019 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3020 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3021 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3022 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3023 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3024 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3025 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3026 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3027 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3028 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3029 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3030 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3031 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3032 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3033 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3034 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3035 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3036 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3037 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3038 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3039 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3040 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3041 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3042 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3043 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3044 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3045 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3046 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3047 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3048 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3049 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3050 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3051 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3052 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3053 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3054 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3055 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3056 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3057 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3058 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3059 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3060 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3061 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3062 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3063 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3064 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3065 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3066 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3067 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3068 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3069 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3070 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3071 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3072 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3073 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3074 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3075 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3076 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3077 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3078 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3079 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3080 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3081 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3082 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3083 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3084 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3085 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3086 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3087 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3088 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3089 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3090 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3091 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3092 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3093 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3094 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3095 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3096 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3097 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3098 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3099 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3100 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3101 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3102 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3103 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3104 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3105 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3106 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3107 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3108 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3109 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3110 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3111 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3112 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3113 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3114 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3115 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3116 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3117 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3118 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3119 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3120 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3121 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3122 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3123 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3124 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3125 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3126 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3127 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3128 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3129 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3130 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3131 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3132 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3133 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3134 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3135 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3136 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3137 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3138 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3139 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3140 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3141 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3142 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3143 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3144 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3145 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3146 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3147 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3148 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3149 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3150 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3151 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3152 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3153 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3154 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3155 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3156 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3157 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3158 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3159 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3160 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3161 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3162 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3163 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3164 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3165 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3166 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3167 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3168 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3169 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3170 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3171 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3172 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3173 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3174 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3175 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3176 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3177 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3178 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3179 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3180 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3181 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3182 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3183 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3184 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3185 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3186 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3187 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3188 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3189 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3190 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3191 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3192 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3193 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3194 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3195 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3196 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3197 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3198 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3199 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3200 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3201 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3202 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3203 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3204 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3205 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3206 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3207 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3208 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3209 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3210 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3211 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3212 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3213 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3214 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3215 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3216 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3217 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3218 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3219 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3220 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3221 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3222 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3223 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3224 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3225 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3226 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3227 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3228 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3229 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3230 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3231 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3232 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3233 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3234 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3235 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3236 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3237 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3238 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3239 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3240 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3241 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3242 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3243 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3244 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3245 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3246 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3247 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3248 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3249 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3250 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3251 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3252 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3253 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3254 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3255 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3256 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3257 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3258 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3259 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3260 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3261 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3262 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3263 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3264 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3265 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3266 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3267 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3268 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3269 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3270 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3271 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3272 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3273 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3274 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3275 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3276 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3277 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3278 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3279 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3280 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3281 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3282 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3283 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3284 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3285 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3286 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3287 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3288 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3289 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3290 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3291 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3292 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3293 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3294 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3295 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3296 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3297 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3298 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3299 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3300 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3301 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3302 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3303 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3304 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3305 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3306 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3307 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3308 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3309 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3310 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3311 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3312 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3313 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3314 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3315 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3316 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3317 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3318 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3319 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3320 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3321 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3322 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3323 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3324 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3325 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3326 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3327 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3328 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3329 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3330 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3331 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3332 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3333 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3334 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3335 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3336 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3337 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3338 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3339 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3340 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3341 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3342 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3343 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3344 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3345 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3346 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3347 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3348 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3349 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3350 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3351 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3352 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3353 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3354 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3355 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3356 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3357 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3358 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3359 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3360 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3361 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3362 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3363 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3364 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3365 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3366 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3367 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3368 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3369 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3370 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3371 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3372 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3373 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3374 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3375 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3376 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3377 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3378 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3379 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3380 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3381 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3382 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3383 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3384 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3385 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3386 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3387 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3388 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3389 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3390 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3391 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3392 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3393 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3394 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3395 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3396 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3397 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3398 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3399 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3400 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3401 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3402 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3403 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3404 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3405 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3406 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3407 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3408 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3409 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3410 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3411 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3412 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3413 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3414 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3415 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3416 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3417 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3418 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3419 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3420 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3421 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3422 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3423 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3424 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3425 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3426 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3427 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3428 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3429 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3430 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3431 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3432 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3433 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3434 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3435 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3436 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3437 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3438 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3439 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3440 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3441 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3442 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3443 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3444 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3445 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3446 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3447 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3448 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3449 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3450 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3451 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3452 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3453 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3454 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3455 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3456 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3457 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3458 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3459 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3460 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3461 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3462 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3463 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3464 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3465 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3466 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3467 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3468 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3469 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3470 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3471 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3472 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3473 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3474 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3475 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3476 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3477 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3478 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3479 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3480 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3481 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3482 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3483 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3484 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3485 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3486 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3487 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3488 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3489 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3490 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3491 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3492 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3493 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3494 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3495 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3496 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3497 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3498 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3499 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3500 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3501 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3502 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3503 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3504 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3505 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3506 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3507 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3508 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3509 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3510 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3511 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3512 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3513 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3514 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3515 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3516 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3517 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3518 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3519 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3520 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3521 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3522 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3523 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3524 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3525 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3526 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3527 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3528 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3529 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3530 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3531 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3532 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3533 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3534 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3535 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3536 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3537 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3538 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3539 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3540 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3541 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3542 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3543 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3544 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3545 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3546 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3547 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3548 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3549 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3550 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3551 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3552 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3553 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3554 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3555 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3556 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3557 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3558 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3559 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3560 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3561 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3562 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3563 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3564 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3565 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3566 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3567 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3568 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3569 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3570 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3571 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3572 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3573 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3574 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3575 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3576 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3577 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3578 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3579 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3580 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3581 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3582 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3583 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3584 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3585 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3586 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3587 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3588 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3589 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3590 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3591 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3592 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3593 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3594 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3595 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3596 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3597 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3598 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3599 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3600 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3601 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3602 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3603 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3604 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3605 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3606 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3607 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3608 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3609 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3610 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3611 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3612 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3613 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3614 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3615 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3616 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3617 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3618 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3619 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3620 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3621 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3622 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3623 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3624 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3625 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3626 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3627 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3628 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3629 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3630 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3631 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3632 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3633 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3634 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3635 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3636 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3637 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3638 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3639 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3640 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3641 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3642 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3643 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3644 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3645 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3646 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3647 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3648 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3649 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3650 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3651 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3652 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3653 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3654 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3655 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3656 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3657 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3658 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3659 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3660 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3661 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3662 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3663 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3664 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3665 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3666 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3667 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3668 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3669 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3670 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3671 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3672 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3673 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3674 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3675 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3676 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3677 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3678 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3679 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3680 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3681 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3682 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3683 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3684 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3685 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3686 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3687 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3688 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3689 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3690 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3691 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3692 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3693 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3694 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3695 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3696 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3697 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3698 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3699 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3700 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3701 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3702 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3703 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3704 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3705 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3706 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3707 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3708 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3709 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3710 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3711 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3712 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3713 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3714 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3715 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3716 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3717 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3718 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3719 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3720 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3721 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3722 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3723 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3724 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3725 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3726 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3727 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3728 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3729 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3730 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3731 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3732 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3733 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3734 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3735 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3736 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3737 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3738 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3739 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3740 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3741 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3742 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3743 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3744 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3745 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3746 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3747 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3748 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3749 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3750 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3751 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3752 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3753 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3754 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3755 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3756 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3757 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3758 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3759 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3760 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3761 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3762 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3763 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3764 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3765 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3766 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3767 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3768 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3769 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3770 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3771 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3772 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3773 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3774 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3775 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3776 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3777 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3778 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3779 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3780 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3781 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3782 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3783 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3784 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3785 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3786 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3787 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3788 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3789 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3790 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3791 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3792 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3793 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3794 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3795 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3796 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3797 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3798 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3799 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3800 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3801 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3802 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3803 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3804 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3805 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3806 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3807 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3808 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3809 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3810 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3811 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3812 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3813 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3814 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3815 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3816 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3817 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3818 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3819 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3820 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3821 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3822 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3823 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3824 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3825 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3826 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3827 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3828 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3829 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3830 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3831 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3832 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3833 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3834 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3835 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3836 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3837 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3838 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3839 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3840 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3841 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3842 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3843 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3844 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3845 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3846 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3847 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3848 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3849 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3850 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3851 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3852 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3853 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3854 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3855 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3856 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3857 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3858 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3859 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3860 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3861 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3862 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3863 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3864 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3865 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3866 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3867 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3868 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3869 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3870 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3871 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3872 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3873 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3874 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3875 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3876 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3877 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3878 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3879 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3880 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3881 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3882 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3883 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3884 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3885 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3886 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3887 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3888 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3889 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3890 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3891 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3892 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3893 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3894 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3895 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3896 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3897 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3898 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3899 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3900 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3901 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3902 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3903 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3904 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3905 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3906 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3907 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3908 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3909 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3910 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3911 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3912 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3913 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3914 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3915 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3916 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3917 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3918 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3919 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3920 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3921 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3922 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3923 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3924 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3925 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3926 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3927 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3928 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3929 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3930 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3931 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3932 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3933 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3934 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3935 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3936 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3937 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3938 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3939 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3940 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3941 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3942 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3943 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3944 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3945 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3946 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3947 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3948 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3949 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3950 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3951 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3952 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3953 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3954 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3955 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3956 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3957 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3958 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3959 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3960 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3961 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3962 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3963 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3964 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3965 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3966 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3967 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3968 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3969 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3970 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3971 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3972 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3973 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3974 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3975 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3976 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3977 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3978 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3979 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3980 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3981 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3982 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3983 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3984 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3985 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3986 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3987 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3988 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3989 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3990 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3991 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3992 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3993 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3994 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3995 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3996 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3997 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3998 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		3999 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4000 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4001 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4002 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4003 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4004 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4005 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4006 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4007 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4008 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4009 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4010 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4011 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4012 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4013 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4014 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4015 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4016 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4017 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4018 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4019 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4020 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4021 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4022 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4023 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4024 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4025 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4026 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4027 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4028 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4029 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4030 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4031 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4032 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4033 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4034 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4035 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4036 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4037 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4038 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4039 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4040 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4041 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4042 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4043 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4044 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4045 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4046 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4047 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4048 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4049 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4050 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4051 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4052 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4053 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4054 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4055 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4056 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4057 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4058 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4059 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4060 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4061 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4062 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4063 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4064 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4065 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4066 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4067 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4068 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4069 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4070 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4071 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4072 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4073 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4074 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4075 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4076 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4077 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4078 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4079 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4080 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4081 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4082 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4083 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4084 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4085 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4086 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4087 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4088 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4089 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4090 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4091 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4092 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4093 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4094 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4095 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4096 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4097 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4098 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4099 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4100 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4101 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4102 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4103 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4104 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4105 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4106 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4107 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4108 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4109 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4110 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4111 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4112 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4113 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4114 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4115 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4116 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4117 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4118 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4119 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4120 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4121 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4122 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4123 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4124 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4125 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4126 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4127 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4128 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4129 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4130 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4131 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4132 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4133 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4134 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4135 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4136 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4137 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4138 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4139 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4140 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4141 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4142 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4143 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4144 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4145 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4146 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4147 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4148 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4149 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4150 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4151 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4152 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4153 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4154 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4155 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4156 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4157 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4158 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4159 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4160 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4161 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4162 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4163 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4164 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4165 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4166 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4167 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4168 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4169 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4170 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4171 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4172 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4173 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4174 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4175 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4176 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4177 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4178 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4179 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4180 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4181 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4182 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4183 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4184 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4185 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4186 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4187 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4188 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4189 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4190 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4191 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4192 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4193 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4194 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4195 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4196 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4197 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4198 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4199 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4200 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4201 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4202 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4203 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4204 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4205 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4206 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4207 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4208 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4209 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4210 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4211 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4212 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4213 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4214 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4215 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4216 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4217 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4218 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4219 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4220 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4221 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4222 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4223 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4224 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4225 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4226 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4227 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4228 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4229 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4230 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4231 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4232 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4233 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4234 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4235 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4236 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4237 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4238 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4239 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4240 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4241 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4242 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4243 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4244 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4245 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4246 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4247 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4248 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4249 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4250 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4251 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4252 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4253 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4254 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4255 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4256 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4257 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4258 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4259 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4260 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4261 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4262 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4263 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4264 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4265 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4266 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4267 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4268 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4269 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4270 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4271 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4272 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4273 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4274 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4275 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4276 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4277 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4278 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4279 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4280 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4281 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4282 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4283 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4284 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4285 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4286 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4287 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4288 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4289 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4290 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4291 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4292 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4293 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4294 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4295 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4296 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4297 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4298 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4299 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4300 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4301 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4302 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4303 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4304 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4305 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4306 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4307 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4308 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4309 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4310 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4311 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4312 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4313 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4314 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4315 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4316 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4317 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4318 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4319 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4320 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4321 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4322 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4323 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4324 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4325 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4326 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4327 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4328 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4329 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4330 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4331 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4332 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4333 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4334 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4335 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4336 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4337 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4338 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4339 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4340 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4341 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4342 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4343 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4344 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4345 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4346 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4347 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4348 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4349 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4350 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4351 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4352 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4353 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4354 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4355 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4356 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4357 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4358 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4359 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4360 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4361 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4362 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4363 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4364 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4365 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4366 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4367 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4368 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4369 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4370 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4371 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4372 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4373 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4374 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4375 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4376 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4377 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4378 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4379 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4380 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4381 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4382 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4383 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4384 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4385 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4386 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4387 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4388 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4389 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4390 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4391 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4392 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4393 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4394 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4395 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4396 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4397 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4398 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4399 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4400 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4401 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4402 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4403 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4404 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4405 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4406 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4407 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4408 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4409 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4410 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4411 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4412 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4413 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4414 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4415 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4416 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4417 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4418 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4419 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4420 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4421 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4422 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4423 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4424 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4425 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4426 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4427 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4428 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4429 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4430 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4431 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4432 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4433 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4434 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4435 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4436 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4437 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4438 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4439 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4440 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4441 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4442 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4443 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4444 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4445 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4446 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4447 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4448 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4449 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4450 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4451 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4452 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4453 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4454 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4455 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4456 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4457 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4458 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4459 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4460 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4461 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4462 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4463 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4464 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4465 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4466 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4467 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4468 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4469 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4470 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4471 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4472 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4473 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4474 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4475 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4476 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4477 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4478 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4479 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4480 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4481 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4482 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4483 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4484 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4485 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4486 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4487 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4488 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4489 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4490 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4491 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4492 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4493 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4494 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4495 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4496 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4497 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4498 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4499 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4500 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4501 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4502 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4503 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4504 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4505 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4506 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4507 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4508 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4509 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4510 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4511 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4512 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4513 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4514 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4515 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4516 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4517 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4518 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4519 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4520 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4521 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4522 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4523 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4524 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4525 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4526 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4527 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4528 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4529 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4530 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4531 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4532 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4533 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4534 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4535 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4536 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4537 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4538 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4539 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4540 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4541 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4542 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4543 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4544 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4545 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4546 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4547 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4548 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4549 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4550 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4551 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4552 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4553 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4554 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4555 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4556 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4557 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4558 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4559 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4560 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4561 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4562 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4563 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4564 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4565 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4566 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4567 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4568 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4569 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4570 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4571 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4572 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4573 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4574 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4575 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4576 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4577 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4578 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4579 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4580 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4581 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4582 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4583 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4584 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4585 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4586 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4587 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4588 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4589 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4590 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4591 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4592 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4593 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4594 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4595 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4596 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4597 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4598 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4599 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4600 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4601 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4602 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4603 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4604 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4605 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4606 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4607 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4608 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4609 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4610 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4611 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4612 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4613 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4614 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4615 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4616 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4617 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4618 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4619 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4620 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4621 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4622 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4623 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4624 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4625 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4626 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4627 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4628 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4629 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4630 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4631 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4632 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4633 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4634 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4635 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4636 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4637 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4638 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4639 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4640 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4641 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4642 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4643 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4644 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4645 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4646 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4647 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4648 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4649 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4650 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4651 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4652 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4653 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4654 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4655 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4656 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4657 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4658 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4659 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4660 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4661 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4662 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4663 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4664 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4665 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4666 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4667 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4668 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4669 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4670 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4671 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4672 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4673 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4674 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4675 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4676 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4677 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4678 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4679 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4680 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4681 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4682 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4683 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4684 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4685 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4686 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4687 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4688 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4689 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4690 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4691 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4692 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4693 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4694 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4695 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4696 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4697 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4698 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4699 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4700 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4701 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4702 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4703 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4704 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4705 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4706 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4707 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4708 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4709 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4710 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4711 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4712 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4713 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4714 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4715 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4716 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4717 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4718 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4719 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4720 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4721 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4722 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4723 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4724 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4725 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4726 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4727 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4728 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4729 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4730 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4731 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4732 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4733 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4734 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4735 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4736 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4737 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4738 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4739 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4740 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4741 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4742 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4743 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4744 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4745 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4746 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4747 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4748 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4749 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4750 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4751 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4752 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4753 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4754 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4755 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4756 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4757 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4758 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4759 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4760 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4761 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4762 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4763 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4764 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4765 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4766 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4767 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4768 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4769 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4770 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4771 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4772 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4773 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4774 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4775 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4776 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4777 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4778 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4779 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4780 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4781 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4782 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4783 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4784 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4785 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4786 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4787 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4788 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4789 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4790 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4791 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4792 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4793 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4794 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4795 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4796 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4797 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4798 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4799 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4800 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4801 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4802 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4803 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4804 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4805 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4806 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4807 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4808 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4809 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4810 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4811 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4812 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4813 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4814 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4815 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4816 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4817 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4818 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4819 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4820 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4821 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4822 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4823 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4824 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4825 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4826 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4827 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4828 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4829 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4830 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4831 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4832 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4833 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4834 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4835 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4836 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4837 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4838 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4839 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4840 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4841 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4842 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4843 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4844 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4845 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4846 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4847 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4848 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4849 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4850 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4851 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4852 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4853 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4854 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4855 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4856 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4857 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4858 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4859 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4860 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4861 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4862 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4863 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4864 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4865 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4866 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4867 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4868 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4869 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4870 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4871 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4872 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4873 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4874 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4875 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4876 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4877 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4878 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4879 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4880 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4881 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4882 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4883 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4884 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4885 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4886 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4887 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4888 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4889 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4890 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4891 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4892 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4893 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4894 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4895 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4896 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4897 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4898 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4899 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4900 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4901 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4902 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4903 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4904 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4905 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4906 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4907 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4908 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4909 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4910 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4911 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4912 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4913 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4914 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4915 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4916 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4917 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4918 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4919 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4920 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4921 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4922 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4923 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4924 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4925 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4926 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4927 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4928 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4929 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4930 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4931 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4932 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4933 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4934 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4935 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4936 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4937 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4938 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4939 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4940 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4941 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4942 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4943 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4944 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4945 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4946 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4947 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4948 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4949 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4950 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4951 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4952 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4953 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4954 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4955 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4956 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4957 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4958 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4959 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4960 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4961 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4962 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4963 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4964 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4965 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4966 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4967 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4968 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4969 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4970 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4971 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4972 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4973 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4974 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4975 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4976 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4977 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4978 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4979 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4980 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4981 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4982 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4983 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4984 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4985 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4986 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4987 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4988 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4989 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4990 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4991 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4992 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4993 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4994 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4995 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4996 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4997 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4998 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		4999 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5000 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5001 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5002 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5003 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5004 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5005 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5006 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5007 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5008 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5009 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5010 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5011 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5012 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5013 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5014 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5015 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5016 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5017 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5018 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5019 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5020 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5021 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5022 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5023 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5024 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5025 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5026 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5027 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5028 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5029 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5030 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5031 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5032 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5033 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5034 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5035 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5036 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5037 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5038 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5039 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5040 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5041 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5042 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5043 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5044 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5045 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5046 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5047 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5048 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5049 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5050 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5051 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5052 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5053 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5054 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5055 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5056 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5057 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5058 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5059 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5060 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5061 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5062 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5063 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5064 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5065 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5066 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5067 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5068 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5069 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5070 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5071 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5072 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5073 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5074 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5075 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5076 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5077 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5078 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5079 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5080 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5081 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5082 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5083 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5084 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5085 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5086 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5087 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5088 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5089 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5090 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5091 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5092 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5093 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5094 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5095 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5096 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5097 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5098 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5099 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5100 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5101 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5102 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5103 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5104 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5105 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5106 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5107 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5108 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5109 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5110 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5111 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5112 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5113 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5114 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5115 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5116 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5117 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5118 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5119 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5120 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5121 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5122 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5123 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5124 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5125 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5126 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5127 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5128 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5129 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5130 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5131 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5132 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5133 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5134 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5135 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5136 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5137 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5138 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5139 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5140 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5141 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5142 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5143 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5144 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5145 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5146 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5147 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5148 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5149 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5150 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5151 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5152 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5153 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5154 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5155 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5156 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5157 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5158 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5159 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5160 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5161 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5162 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5163 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5164 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5165 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5166 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5167 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5168 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5169 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5170 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5171 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5172 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5173 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5174 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5175 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5176 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5177 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5178 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5179 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5180 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5181 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5182 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5183 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5184 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5185 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5186 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5187 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5188 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5189 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5190 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5191 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5192 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5193 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5194 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5195 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5196 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5197 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5198 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5199 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5200 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5201 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5202 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5203 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5204 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5205 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5206 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5207 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5208 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5209 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5210 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5211 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5212 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5213 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5214 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5215 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5216 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5217 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5218 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5219 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5220 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5221 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5222 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5223 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5224 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5225 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5226 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5227 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5228 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5229 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5230 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5231 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5232 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5233 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5234 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5235 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5236 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5237 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5238 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5239 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5240 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5241 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5242 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5243 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5244 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5245 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5246 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5247 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5248 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5249 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5250 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5251 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5252 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5253 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5254 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5255 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5256 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5257 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5258 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5259 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5260 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5261 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5262 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5263 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5264 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5265 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5266 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5267 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5268 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5269 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5270 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5271 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5272 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5273 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5274 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5275 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5276 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5277 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5278 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5279 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5280 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5281 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5282 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5283 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5284 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5285 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5286 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5287 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5288 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5289 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5290 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5291 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5292 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5293 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5294 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5295 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5296 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5297 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5298 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5299 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5300 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5301 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5302 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5303 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5304 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5305 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5306 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5307 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5308 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5309 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5310 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5311 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5312 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5313 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5314 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5315 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5316 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5317 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5318 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5319 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5320 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5321 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5322 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5323 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5324 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5325 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5326 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5327 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5328 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5329 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5330 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5331 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5332 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5333 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5334 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5335 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5336 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5337 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5338 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5339 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5340 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5341 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5342 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5343 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5344 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5345 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5346 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5347 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5348 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5349 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5350 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5351 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5352 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5353 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5354 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5355 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5356 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5357 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5358 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5359 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5360 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5361 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5362 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5363 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5364 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5365 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5366 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5367 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5368 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5369 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5370 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5371 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5372 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5373 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5374 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5375 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5376 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5377 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5378 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5379 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5380 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5381 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5382 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5383 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5384 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5385 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5386 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5387 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5388 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5389 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5390 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5391 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5392 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5393 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5394 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5395 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5396 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5397 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5398 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5399 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5400 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5401 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5402 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5403 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5404 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5405 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5406 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5407 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5408 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5409 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5410 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5411 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5412 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5413 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5414 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5415 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5416 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5417 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5418 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5419 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5420 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5421 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5422 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5423 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5424 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5425 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5426 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5427 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5428 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5429 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5430 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5431 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5432 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5433 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5434 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5435 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5436 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5437 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5438 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5439 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5440 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5441 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5442 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5443 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5444 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5445 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5446 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5447 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5448 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5449 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5450 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5451 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5452 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5453 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5454 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5455 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5456 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5457 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5458 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5459 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5460 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5461 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5462 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5463 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5464 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5465 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5466 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5467 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5468 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5469 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5470 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5471 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5472 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5473 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5474 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5475 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5476 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5477 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5478 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5479 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5480 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5481 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5482 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5483 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5484 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5485 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5486 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5487 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5488 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5489 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5490 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5491 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5492 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5493 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5494 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5495 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5496 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5497 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5498 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5499 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5500 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5501 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5502 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5503 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5504 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5505 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5506 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5507 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5508 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5509 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5510 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5511 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5512 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5513 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5514 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5515 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5516 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5517 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5518 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5519 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5520 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5521 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5522 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5523 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5524 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5525 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5526 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5527 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5528 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5529 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5530 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5531 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5532 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5533 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5534 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5535 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5536 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5537 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5538 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5539 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5540 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5541 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5542 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5543 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5544 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5545 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5546 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5547 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5548 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5549 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5550 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5551 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5552 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5553 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5554 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5555 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5556 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5557 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5558 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5559 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5560 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5561 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5562 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5563 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5564 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5565 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5566 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5567 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5568 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5569 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5570 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5571 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5572 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5573 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5574 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5575 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5576 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5577 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5578 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5579 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5580 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5581 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5582 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5583 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5584 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5585 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5586 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5587 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5588 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5589 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5590 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5591 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5592 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5593 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5594 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5595 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5596 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5597 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5598 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5599 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5600 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5601 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5602 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5603 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5604 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5605 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5606 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5607 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5608 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5609 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5610 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5611 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5612 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5613 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5614 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5615 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5616 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5617 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5618 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5619 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5620 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5621 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5622 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5623 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5624 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5625 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5626 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5627 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5628 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5629 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5630 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5631 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5632 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5633 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5634 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5635 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5636 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5637 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5638 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5639 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5640 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5641 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5642 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5643 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5644 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5645 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5646 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5647 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5648 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5649 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5650 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5651 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5652 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5653 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5654 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5655 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5656 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5657 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5658 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5659 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5660 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5661 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5662 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5663 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5664 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5665 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5666 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5667 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5668 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5669 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5670 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5671 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5672 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5673 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5674 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5675 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5676 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5677 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5678 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5679 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5680 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5681 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5682 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5683 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5684 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5685 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5686 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5687 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5688 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5689 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5690 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5691 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5692 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5693 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5694 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5695 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5696 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5697 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5698 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5699 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5700 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5701 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5702 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5703 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5704 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5705 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5706 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5707 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5708 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5709 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5710 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5711 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5712 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5713 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5714 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5715 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5716 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5717 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5718 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5719 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5720 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5721 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5722 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5723 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5724 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5725 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5726 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5727 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5728 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5729 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5730 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5731 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5732 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5733 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5734 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5735 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5736 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5737 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5738 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5739 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5740 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5741 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5742 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5743 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5744 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5745 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5746 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5747 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5748 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5749 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5750 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5751 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5752 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5753 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5754 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5755 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5756 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5757 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5758 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5759 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5760 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5761 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5762 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5763 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5764 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5765 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5766 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5767 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5768 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5769 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5770 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5771 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5772 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5773 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5774 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5775 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5776 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5777 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5778 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5779 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5780 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5781 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5782 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5783 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5784 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5785 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5786 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5787 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5788 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5789 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5790 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5791 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5792 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5793 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5794 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5795 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5796 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5797 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5798 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5799 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5800 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5801 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5802 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5803 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5804 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5805 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5806 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5807 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5808 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5809 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5810 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5811 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5812 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5813 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5814 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5815 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5816 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5817 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5818 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5819 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5820 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5821 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5822 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5823 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5824 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5825 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5826 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5827 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5828 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5829 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5830 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5831 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5832 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5833 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5834 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5835 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5836 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5837 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5838 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5839 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5840 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5841 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5842 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5843 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5844 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5845 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5846 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5847 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5848 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5849 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5850 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5851 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5852 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5853 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5854 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5855 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5856 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5857 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5858 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5859 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5860 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5861 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5862 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5863 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5864 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5865 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5866 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5867 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5868 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5869 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5870 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5871 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5872 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5873 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5874 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5875 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5876 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5877 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5878 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5879 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5880 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5881 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5882 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5883 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5884 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5885 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5886 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5887 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5888 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5889 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5890 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5891 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5892 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5893 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5894 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5895 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5896 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5897 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5898 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5899 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5900 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5901 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5902 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5903 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5904 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5905 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5906 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5907 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5908 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5909 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5910 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5911 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5912 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5913 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5914 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5915 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5916 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5917 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5918 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5919 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5920 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5921 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5922 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5923 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5924 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5925 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5926 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5927 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5928 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5929 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5930 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5931 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5932 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5933 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5934 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5935 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5936 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5937 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5938 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5939 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5940 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5941 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5942 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5943 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5944 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5945 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5946 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5947 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5948 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5949 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5950 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5951 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5952 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5953 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5954 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5955 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5956 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5957 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5958 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5959 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5960 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5961 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5962 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5963 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5964 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5965 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5966 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5967 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5968 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5969 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5970 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5971 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5972 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5973 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5974 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5975 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5976 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5977 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5978 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5979 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5980 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5981 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5982 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5983 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5984 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5985 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5986 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5987 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5988 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5989 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5990 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5991 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5992 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5993 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5994 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5995 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5996 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5997 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5998 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		5999 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6000 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6001 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6002 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6003 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6004 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6005 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6006 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6007 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6008 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6009 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6010 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6011 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6012 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6013 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6014 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6015 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6016 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6017 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6018 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6019 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6020 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6021 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6022 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6023 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6024 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6025 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6026 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6027 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6028 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6029 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6030 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6031 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6032 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6033 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6034 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6035 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6036 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6037 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6038 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6039 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6040 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6041 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6042 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6043 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6044 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6045 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6046 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6047 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6048 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6049 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6050 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6051 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6052 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6053 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6054 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6055 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6056 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6057 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6058 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6059 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6060 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6061 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6062 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6063 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6064 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6065 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6066 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6067 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6068 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6069 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6070 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6071 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6072 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6073 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6074 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6075 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6076 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6077 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6078 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6079 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6080 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6081 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6082 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6083 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6084 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6085 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6086 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6087 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6088 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6089 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6090 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6091 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6092 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6093 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6094 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6095 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6096 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6097 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6098 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6099 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6100 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6101 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6102 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6103 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6104 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6105 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6106 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6107 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6108 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6109 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6110 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6111 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6112 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6113 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6114 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6115 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6116 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6117 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6118 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6119 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6120 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6121 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6122 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6123 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6124 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6125 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6126 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6127 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6128 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6129 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6130 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6131 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6132 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6133 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6134 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6135 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6136 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6137 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6138 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6139 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6140 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6141 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6142 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6143 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6144 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6145 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6146 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6147 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6148 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6149 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6150 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6151 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6152 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6153 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6154 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6155 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6156 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6157 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6158 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6159 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6160 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6161 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6162 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6163 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6164 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6165 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6166 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6167 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6168 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6169 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6170 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6171 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6172 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6173 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6174 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6175 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6176 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6177 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6178 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6179 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6180 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6181 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6182 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6183 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6184 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6185 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6186 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6187 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6188 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6189 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6190 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6191 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6192 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6193 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6194 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6195 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6196 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6197 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6198 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6199 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6200 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6201 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6202 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6203 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6204 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6205 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6206 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		6207 =>	"00000000000000000000000000000000", -- z: 0 rot: 0 ptr: 0
		others => "00000000000000000000000000000000"
	);

begin

	process( clk_i ) begin
		if rising_edge( clk_i ) then
--			if we_i = '1' then
--				mem( to_integer( unsigned( addr_i ) ) ) <= data_o;
--			else
				data_o <= mem( to_integer( unsigned( addr_i ) ) );
--			end if;
		end if; 
	end process;

end architecture arch;